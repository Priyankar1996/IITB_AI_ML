-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity readModule1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    index : in  std_logic_vector(7 downto 0);
    address : in  std_logic_vector(31 downto 0);
    data : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(14 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readModule1;
architecture readModule1_arch of readModule1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 40)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  -- output port buffer signals
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  signal readModule1_CP_26_start: Boolean;
  signal readModule1_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_28_index_0_scale_req_0 : boolean;
  signal array_obj_ref_28_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_28_index_0_scale_req_1 : boolean;
  signal array_obj_ref_28_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_28_index_sum_1_req_0 : boolean;
  signal array_obj_ref_28_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_28_index_sum_1_req_1 : boolean;
  signal array_obj_ref_28_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_28_index_offset_req_0 : boolean;
  signal array_obj_ref_28_index_offset_ack_0 : boolean;
  signal array_obj_ref_28_index_offset_req_1 : boolean;
  signal array_obj_ref_28_index_offset_ack_1 : boolean;
  signal addr_of_29_final_reg_req_0 : boolean;
  signal addr_of_29_final_reg_ack_0 : boolean;
  signal addr_of_29_final_reg_req_1 : boolean;
  signal addr_of_29_final_reg_ack_1 : boolean;
  signal ptr_deref_33_load_0_req_0 : boolean;
  signal ptr_deref_33_load_0_ack_0 : boolean;
  signal ptr_deref_33_load_0_req_1 : boolean;
  signal ptr_deref_33_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readModule1_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 40) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= index;
  index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= address;
  address_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(tag_length + 39 downto 40) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 39 downto 40);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 3) := (0 => 8,1 => 8,2 => 1,3 => 8);
    constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 8);
    constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 4); -- 
  begin -- 
    preds <= index_update_enable & address_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readModule1_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readModule1_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= data_buffer;
  data <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule1_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  data_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "data_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_data_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => data_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 8,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readModule1_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule1_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readModule1_CP_26: Block -- control-path 
    signal readModule1_CP_26_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    readModule1_CP_26_elements(0) <= readModule1_CP_26_start;
    readModule1_CP_26_symbol <= readModule1_CP_26_elements(30);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	13 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	6 
    -- CP-element group 1: 	17 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resized_2
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scaled_2
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_computed_2
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/$entry
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resized_0
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_computed_0
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resize_2/$entry
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resize_2/$exit
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resize_2/index_resize_req
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_resize_2/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_2/$entry
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_2/$exit
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_2/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_2/scale_rename_ack
      -- 
    readModule1_CP_26_elements(1) <= readModule1_CP_26_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	27 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_30_to_assign_stmt_34/index_update_enable
      -- CP-element group 2: 	 assign_stmt_30_to_assign_stmt_34/index_update_enable_out
      -- 
    readModule1_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readModule1_CP_26_elements(8);
      gj_readModule1_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	15 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	28 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_30_to_assign_stmt_34/address_update_enable
      -- CP-element group 3: 	 assign_stmt_30_to_assign_stmt_34/address_update_enable_out
      -- 
    readModule1_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readModule1_CP_26_elements(15);
      gj_readModule1_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	29 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	23 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_30_to_assign_stmt_34/data_update_enable
      -- CP-element group 4: 	 assign_stmt_30_to_assign_stmt_34/data_update_enable_in
      -- 
    readModule1_CP_26_elements(4) <= readModule1_CP_26_elements(29);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	20 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	20 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_sample_start_
      -- CP-element group 5: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_request/$entry
      -- CP-element group 5: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_request/req
      -- 
    req_113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(5), ack => addr_of_29_final_reg_req_0); -- 
    readModule1_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(7) & readModule1_CP_26_elements(20);
      gj_readModule1_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	21 
    -- CP-element group 6: 	24 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_update_start_
      -- CP-element group 6: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_complete/$entry
      -- CP-element group 6: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_complete/req
      -- 
    req_118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(6), ack => addr_of_29_final_reg_req_1); -- 
    readModule1_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(1) & readModule1_CP_26_elements(21) & readModule1_CP_26_elements(24);
      gj_readModule1_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	16 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	17 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_root_address_calculated
      -- CP-element group 7: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_offset_calculated
      -- CP-element group 7: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_base_plus_offset/$entry
      -- CP-element group 7: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_base_plus_offset/$exit
      -- CP-element group 7: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_base_plus_offset/sum_rename_req
      -- CP-element group 7: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_base_plus_offset/sum_rename_ack
      -- 
    readModule1_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 8);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(19) & readModule1_CP_26_elements(16);
      gj_readModule1_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	15 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scaled_0
      -- 
    readModule1_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(12) & readModule1_CP_26_elements(15);
      gj_readModule1_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_sample_start
      -- CP-element group 9: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_Sample/rr
      -- 
    rr_59_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_59_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(9), ack => array_obj_ref_28_index_0_scale_req_0); -- 
    readModule1_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(1) & readModule1_CP_26_elements(11);
      gj_readModule1_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_update_start
      -- CP-element group 10: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_Update/$entry
      -- CP-element group 10: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_Update/cr
      -- 
    cr_64_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_64_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(10), ack => array_obj_ref_28_index_0_scale_req_1); -- 
    readModule1_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(1) & readModule1_CP_26_elements(12);
      gj_readModule1_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	26 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_sample_complete
      -- CP-element group 11: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_Sample/ra
      -- 
    ra_60_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_28_index_0_scale_ack_0, ack => readModule1_CP_26_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_update_complete
      -- CP-element group 12: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_Update/$exit
      -- CP-element group 12: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_index_scale_0_Update/ca
      -- 
    ca_65_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_28_index_0_scale_ack_1, ack => readModule1_CP_26_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	1 
    -- CP-element group 13: 	8 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_sample_start
      -- CP-element group 13: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_Sample/rr
      -- 
    rr_86_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_86_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(13), ack => array_obj_ref_28_index_sum_1_req_0); -- 
    readModule1_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(1) & readModule1_CP_26_elements(8) & readModule1_CP_26_elements(15);
      gj_readModule1_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_update_start
      -- CP-element group 14: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_Update/$entry
      -- CP-element group 14: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_Update/cr
      -- 
    cr_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(14), ack => array_obj_ref_28_index_sum_1_req_1); -- 
    readModule1_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(1) & readModule1_CP_26_elements(18) & readModule1_CP_26_elements(16);
      gj_readModule1_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	26 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: 	13 
    -- CP-element group 15: 	8 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_sample_complete
      -- CP-element group 15: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_Sample/$exit
      -- CP-element group 15: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_Sample/ra
      -- 
    ra_87_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_28_index_sum_1_ack_0, ack => readModule1_CP_26_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: 	18 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_update_complete
      -- CP-element group 16: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_Update/$exit
      -- CP-element group 16: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_partial_sum_1_Update/ca
      -- CP-element group 16: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_Sample/$entry
      -- CP-element group 16: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_Sample/req
      -- 
    ca_92_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_28_index_sum_1_ack_1, ack => readModule1_CP_26_elements(16)); -- 
    req_98_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_98_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(16), ack => array_obj_ref_28_index_offset_req_0); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	7 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_update_start
      -- CP-element group 17: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_Update/$entry
      -- CP-element group 17: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_Update/req
      -- 
    req_103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(17), ack => array_obj_ref_28_index_offset_req_1); -- 
    readModule1_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(1) & readModule1_CP_26_elements(7) & readModule1_CP_26_elements(20);
      gj_readModule1_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	26 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_Sample/ack
      -- 
    ack_99_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_28_index_offset_ack_0, ack => readModule1_CP_26_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	7 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 assign_stmt_30_to_assign_stmt_34/array_obj_ref_28_final_index_sum_regn_Update/ack
      -- 
    ack_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_28_index_offset_ack_1, ack => readModule1_CP_26_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	5 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	5 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_sample_completed_
      -- CP-element group 20: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_request/$exit
      -- CP-element group 20: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_request/ack
      -- 
    ack_114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_29_final_reg_ack_0, ack => readModule1_CP_26_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	6 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_update_completed_
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_complete/$exit
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/addr_of_29_complete/ack
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_address_calculated
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_word_address_calculated
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_root_address_calculated
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_address_resized
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_addr_resize/$entry
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_addr_resize/$exit
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_plus_offset/$entry
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_plus_offset/$exit
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_word_addrgen/$entry
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_word_addrgen/$exit
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_word_addrgen/root_register_req
      -- CP-element group 21: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_word_addrgen/root_register_ack
      -- 
    ack_119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_29_final_reg_ack_1, ack => readModule1_CP_26_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_sample_start_
      -- CP-element group 22: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Sample/$entry
      -- CP-element group 22: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Sample/word_access_start/$entry
      -- CP-element group 22: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Sample/word_access_start/word_0/$entry
      -- CP-element group 22: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Sample/word_access_start/word_0/rr
      -- 
    rr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(22), ack => ptr_deref_33_load_0_req_0); -- 
    readModule1_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(21) & readModule1_CP_26_elements(24);
      gj_readModule1_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	4 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_update_start_
      -- CP-element group 23: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/$entry
      -- CP-element group 23: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/word_access_complete/$entry
      -- CP-element group 23: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/word_access_complete/word_0/$entry
      -- CP-element group 23: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/word_access_complete/word_0/cr
      -- 
    cr_163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_26_elements(23), ack => ptr_deref_33_load_0_req_1); -- 
    readModule1_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(4) & readModule1_CP_26_elements(25);
      gj_readModule1_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: 	6 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_sample_completed_
      -- CP-element group 24: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Sample/$exit
      -- CP-element group 24: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Sample/word_access_start/$exit
      -- CP-element group 24: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Sample/word_access_start/word_0/ra
      -- 
    ra_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_33_load_0_ack_0, ack => readModule1_CP_26_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_update_completed_
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/$exit
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/word_access_complete/$exit
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/ptr_deref_33_Merge/$entry
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/ptr_deref_33_Merge/$exit
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/ptr_deref_33_Merge/merge_req
      -- CP-element group 25: 	 assign_stmt_30_to_assign_stmt_34/ptr_deref_33_Update/ptr_deref_33_Merge/merge_ack
      -- 
    ca_164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_33_load_0_ack_1, ack => readModule1_CP_26_elements(25)); -- 
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	11 
    -- CP-element group 26: 	25 
    -- CP-element group 26: 	15 
    -- CP-element group 26: 	18 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	30 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 assign_stmt_30_to_assign_stmt_34/$exit
      -- 
    readModule1_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 8,1 => 8,2 => 8,3 => 8);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= readModule1_CP_26_elements(11) & readModule1_CP_26_elements(25) & readModule1_CP_26_elements(15) & readModule1_CP_26_elements(18);
      gj_readModule1_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_26_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  place  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 index_update_enable
      -- 
    readModule1_CP_26_elements(27) <= readModule1_CP_26_elements(2);
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	3 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 address_update_enable
      -- 
    readModule1_CP_26_elements(28) <= readModule1_CP_26_elements(3);
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	4 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 data_update_enable
      -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	26 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 $exit
      -- 
    readModule1_CP_26_elements(30) <= readModule1_CP_26_elements(26);
    --  hookup: inputs to control-path 
    readModule1_CP_26_elements(29) <= data_update_enable;
    -- hookup: output from control-path 
    index_update_enable <= readModule1_CP_26_elements(27);
    address_update_enable <= readModule1_CP_26_elements(28);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_address_27_resized : std_logic_vector(14 downto 0);
    signal R_address_27_scaled : std_logic_vector(14 downto 0);
    signal array_obj_ref_28_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_28_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_28_index_partial_sum_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_28_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_28_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_28_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_28_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_28_root_address : std_logic_vector(14 downto 0);
    signal ptr_30 : std_logic_vector(31 downto 0);
    signal ptr_deref_33_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_33_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_33_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_33_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_33_word_offset_0 : std_logic_vector(14 downto 0);
    signal type_cast_24_resized : std_logic_vector(14 downto 0);
    signal type_cast_24_scaled : std_logic_vector(14 downto 0);
    signal type_cast_24_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_28_constant_part_of_offset <= "000000000000000";
    array_obj_ref_28_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_28_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_28_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_28_resized_base_address <= "000000000000000";
    ptr_deref_33_word_offset_0 <= "000000000000000";
    addr_of_29_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_29_final_reg_req_0;
      addr_of_29_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_29_final_reg_req_1;
      addr_of_29_final_reg_ack_1<= rack(0);
      addr_of_29_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_29_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_28_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_30,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_24_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := index_buffer(7 downto 0);
      type_cast_24_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_28_index_0_resize
    process(type_cast_24_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_24_wire;
      ov := iv(14 downto 0);
      type_cast_24_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_28_index_2_rename
    process(R_address_27_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_27_resized;
      ov(14 downto 0) := iv;
      R_address_27_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_28_index_2_resize
    process(address_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_buffer;
      ov := iv(14 downto 0);
      R_address_27_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_28_root_address_inst
    process(array_obj_ref_28_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_28_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_28_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_33_addr_0
    process(ptr_deref_33_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_33_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_33_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_33_base_resize
    process(ptr_30) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_30;
      ov := iv(14 downto 0);
      ptr_deref_33_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_33_gather_scatter
    process(ptr_deref_33_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_33_data_0;
      ov(63 downto 0) := iv;
      data_buffer <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_33_root_address_inst
    process(ptr_deref_33_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_33_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_33_root_address <= ov(14 downto 0);
      --
    end process;
    -- shared split operator group (0) : array_obj_ref_28_index_0_scale 
    ApIntMul_group_0: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_24_resized;
      type_cast_24_scaled <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_28_index_0_scale_req_0;
      array_obj_ref_28_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_28_index_0_scale_req_1;
      array_obj_ref_28_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_0_gI: SplitGuardInterface generic map(name => "ApIntMul_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "100000000000000",
          constant_width => 15,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_28_index_offset 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= array_obj_ref_28_index_partial_sum_1;
      array_obj_ref_28_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_28_index_offset_req_0;
      array_obj_ref_28_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_28_index_offset_req_1;
      array_obj_ref_28_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "000000000000000",
          constant_width => 15,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_28_index_sum_1 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_27_scaled & type_cast_24_scaled;
      array_obj_ref_28_index_partial_sum_1 <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_28_index_sum_1_req_0;
      array_obj_ref_28_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_28_index_sum_1_req_1;
      array_obj_ref_28_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 15, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared load operator group (0) : ptr_deref_33_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_33_load_0_req_0;
      ptr_deref_33_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_33_load_0_req_1;
      ptr_deref_33_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_33_word_address_0;
      ptr_deref_33_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 15,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(14 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end readModule1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_173_start: Boolean;
  signal timer_CP_173_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_39_load_0_req_0 : boolean;
  signal LOAD_count_39_load_0_ack_0 : boolean;
  signal LOAD_count_39_load_0_req_1 : boolean;
  signal LOAD_count_39_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_173_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_173_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_173_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_173_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_173: Block -- control-path 
    signal timer_CP_173_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_173_elements(0) <= timer_CP_173_start;
    timer_CP_173_symbol <= timer_CP_173_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_40/$entry
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_sample_start_
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_update_start_
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_Update/$entry
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_40/LOAD_count_39_Update/word_access_complete/word_0/cr
      -- 
    rr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_173_elements(0), ack => LOAD_count_39_load_0_req_0); -- 
    cr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_173_elements(0), ack => LOAD_count_39_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_40/LOAD_count_39_sample_completed_
      -- CP-element group 1: 	 assign_stmt_40/LOAD_count_39_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_40/LOAD_count_39_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_40/LOAD_count_39_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_40/LOAD_count_39_Sample/word_access_start/word_0/ra
      -- 
    ra_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_39_load_0_ack_0, ack => timer_CP_173_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_40/$exit
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_update_completed_
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_Update/$exit
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_Update/LOAD_count_39_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_Update/LOAD_count_39_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_Update/LOAD_count_39_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_40/LOAD_count_39_Update/LOAD_count_39_Merge/merge_ack
      -- 
    ca_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_39_load_0_ack_1, ack => timer_CP_173_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_39_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_39_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_39_word_address_0 <= "0";
    -- equivalence LOAD_count_39_gather_scatter
    process(LOAD_count_39_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_39_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_39_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_39_load_0_req_0;
      LOAD_count_39_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_39_load_0_req_1;
      LOAD_count_39_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_39_word_address_0;
      LOAD_count_39_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_212_start: Boolean;
  signal timerDaemon_CP_212_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_44_branch_req_0 : boolean;
  signal phi_stmt_46_req_1 : boolean;
  signal phi_stmt_46_req_0 : boolean;
  signal phi_stmt_46_ack_0 : boolean;
  signal ADD_u64_u64_52_inst_req_0 : boolean;
  signal ADD_u64_u64_52_inst_ack_0 : boolean;
  signal ADD_u64_u64_52_inst_req_1 : boolean;
  signal ADD_u64_u64_52_inst_ack_1 : boolean;
  signal STORE_count_54_store_0_req_0 : boolean;
  signal STORE_count_54_store_0_ack_0 : boolean;
  signal STORE_count_54_store_0_req_1 : boolean;
  signal STORE_count_54_store_0_ack_1 : boolean;
  signal do_while_stmt_44_branch_ack_0 : boolean;
  signal do_while_stmt_44_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_212_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_212_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_212_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_212_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_212: Block -- control-path 
    signal timerDaemon_CP_212_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_212_elements(0) <= timerDaemon_CP_212_start;
    timerDaemon_CP_212_symbol <= timerDaemon_CP_212_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_43/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/branch_block_stmt_43__entry__
      -- CP-element group 0: 	 branch_block_stmt_43/do_while_stmt_44__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_43/$exit
      -- CP-element group 1: 	 branch_block_stmt_43/branch_block_stmt_43__exit__
      -- CP-element group 1: 	 branch_block_stmt_43/do_while_stmt_44__exit__
      -- 
    timerDaemon_CP_212_elements(1) <= timerDaemon_CP_212_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_43/do_while_stmt_44/$entry
      -- CP-element group 2: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44__entry__
      -- 
    timerDaemon_CP_212_elements(2) <= timerDaemon_CP_212_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44__exit__
      -- 
    -- Element group timerDaemon_CP_212_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_43/do_while_stmt_44/loop_back
      -- 
    -- Element group timerDaemon_CP_212_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	38 
    -- CP-element group 5: 	37 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_43/do_while_stmt_44/condition_done
      -- CP-element group 5: 	 branch_block_stmt_43/do_while_stmt_44/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_43/do_while_stmt_44/loop_taken/$entry
      -- 
    timerDaemon_CP_212_elements(5) <= timerDaemon_CP_212_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_43/do_while_stmt_44/loop_body_done
      -- 
    timerDaemon_CP_212_elements(6) <= timerDaemon_CP_212_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_212_elements(7) <= timerDaemon_CP_212_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_212_elements(8) <= timerDaemon_CP_212_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_212_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	35 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/condition_evaluated
      -- 
    condition_evaluated_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_212_elements(10), ack => do_while_stmt_44_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_212_elements(15) & timerDaemon_CP_212_elements(35);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_212_elements(12) & timerDaemon_CP_212_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_212_elements(9) & timerDaemon_CP_212_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start_
      -- CP-element group 13: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_212_elements(9) & timerDaemon_CP_212_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_212_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_212_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_trigger
      -- 
    timerDaemon_CP_212_elements(16) <= timerDaemon_CP_212_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req_ps
      -- 
    phi_stmt_46_loopback_sample_req_251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_loopback_sample_req_251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_212_elements(17), ack => phi_stmt_46_req_1); -- 
    -- Element group timerDaemon_CP_212_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_trigger
      -- 
    timerDaemon_CP_212_elements(18) <= timerDaemon_CP_212_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req_ps
      -- 
    phi_stmt_46_entry_sample_req_254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_entry_sample_req_254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_212_elements(19), ack => phi_stmt_46_req_0); -- 
    -- Element group timerDaemon_CP_212_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack_ps
      -- 
    phi_stmt_46_phi_mux_ack_257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_46_ack_0, ack => timerDaemon_CP_212_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_completed_
      -- 
    -- Element group timerDaemon_CP_212_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_start_
      -- 
    -- Element group timerDaemon_CP_212_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_completed__ps
      -- 
    timerDaemon_CP_212_elements(23) <= timerDaemon_CP_212_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_completed_
      -- 
    -- Element group timerDaemon_CP_212_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_212_elements(22), ack => timerDaemon_CP_212_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_212_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_update_start__ps
      -- 
    -- Element group timerDaemon_CP_212_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_Sample/rr
      -- 
    rr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_212_elements(27), ack => ADD_u64_u64_52_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_212_elements(25) & timerDaemon_CP_212_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_update_start_
      -- CP-element group 28: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_Update/cr
      -- 
    cr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_212_elements(28), ack => ADD_u64_u64_52_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_212_elements(26) & timerDaemon_CP_212_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_Sample/ra
      -- 
    ra_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_52_inst_ack_0, ack => timerDaemon_CP_212_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/ADD_u64_u64_52_Update/ca
      -- 
    ca_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_52_inst_ack_1, ack => timerDaemon_CP_212_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/STORE_count_54_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/STORE_count_54_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/STORE_count_54_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/STORE_count_54_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/word_access_start/word_0/rr
      -- 
    rr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_212_elements(31), ack => STORE_count_54_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_212_elements(9) & timerDaemon_CP_212_elements(15) & timerDaemon_CP_212_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_update_start_
      -- CP-element group 32: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Update/word_access_complete/word_0/cr
      -- 
    cr_317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_212_elements(32), ack => STORE_count_54_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_212_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Sample/word_access_start/word_0/ra
      -- 
    ra_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_54_store_0_ack_0, ack => timerDaemon_CP_212_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/STORE_count_54_Update/word_access_complete/word_0/ca
      -- 
    ca_318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_54_store_0_ack_1, ack => timerDaemon_CP_212_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_212_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_212_elements(9), ack => timerDaemon_CP_212_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_43/do_while_stmt_44/do_while_stmt_44_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_212_elements(14) & timerDaemon_CP_212_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_212_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_43/do_while_stmt_44/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_43/do_while_stmt_44/loop_exit/ack
      -- 
    ack_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_0, ack => timerDaemon_CP_212_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_43/do_while_stmt_44/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_43/do_while_stmt_44/loop_taken/ack
      -- 
    ack_327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_1, ack => timerDaemon_CP_212_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_43/do_while_stmt_44/$exit
      -- 
    timerDaemon_CP_212_elements(39) <= timerDaemon_CP_212_elements(3);
    timerDaemon_do_while_stmt_44_terminator_328: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_44_terminator_328", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_212_elements(6),loop_continue => timerDaemon_CP_212_elements(38),loop_terminate => timerDaemon_CP_212_elements(37),loop_back => timerDaemon_CP_212_elements(4),loop_exit => timerDaemon_CP_212_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_46_phi_seq_285_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_212_elements(18);
      timerDaemon_CP_212_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_212_elements(21);
      timerDaemon_CP_212_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_212_elements(23);
      timerDaemon_CP_212_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_212_elements(16);
      timerDaemon_CP_212_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_212_elements(29);
      timerDaemon_CP_212_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_212_elements(30);
      timerDaemon_CP_212_elements(17) <= phi_mux_reqs(1);
      phi_stmt_46_phi_seq_285 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_46_phi_seq_285") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_212_elements(11), 
          phi_sample_ack => timerDaemon_CP_212_elements(14), 
          phi_update_req => timerDaemon_CP_212_elements(13), 
          phi_update_ack => timerDaemon_CP_212_elements(15), 
          phi_mux_ack => timerDaemon_CP_212_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_237_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_212_elements(7);
        preds(1)  <= timerDaemon_CP_212_elements(8);
        entry_tmerge_237 : transition_merge -- 
          generic map(name => " entry_tmerge_237")
          port map (preds => preds, symbol_out => timerDaemon_CP_212_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_52_wire : std_logic_vector(63 downto 0);
    signal STORE_count_54_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_54_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_51_wire_constant : std_logic_vector(63 downto 0);
    signal konst_58_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_46 : std_logic_vector(63 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_54_word_address_0 <= "0";
    konst_51_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_58_wire_constant <= "1";
    type_cast_49_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_46: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_49_wire_constant & ADD_u64_u64_52_wire;
      req <= phi_stmt_46_req_0 & phi_stmt_46_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_46",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_46_ack_0,
          idata => idata,
          odata => ncount_46,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_46
    -- equivalence STORE_count_54_gather_scatter
    process(ncount_46) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_46;
      ov(63 downto 0) := iv;
      STORE_count_54_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_44_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_58_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_44_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_44_branch_req_0,
          ack0 => do_while_stmt_44_branch_ack_0,
          ack1 => do_while_stmt_44_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_52_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_46;
      ADD_u64_u64_52_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_52_inst_req_0;
      ADD_u64_u64_52_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_52_inst_req_1;
      ADD_u64_u64_52_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_54_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_54_store_0_req_0;
      STORE_count_54_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_54_store_0_req_1;
      STORE_count_54_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_54_word_address_0;
      data_in <= STORE_count_54_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity writeModule1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    index : in  std_logic_vector(7 downto 0);
    address : in  std_logic_vector(31 downto 0);
    data : in  std_logic_vector(63 downto 0);
    done : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(14 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeModule1;
architecture writeModule1_arch of writeModule1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 104)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  -- output port buffer signals
  signal done_buffer :  std_logic_vector(0 downto 0);
  signal done_update_enable: Boolean;
  signal writeModule1_CP_329_start: Boolean;
  signal writeModule1_CP_329_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal BITSEL_u8_u1_83_inst_req_0 : boolean;
  signal BITSEL_u8_u1_83_inst_ack_0 : boolean;
  signal BITSEL_u8_u1_83_inst_req_1 : boolean;
  signal BITSEL_u8_u1_83_inst_ack_1 : boolean;
  signal array_obj_ref_73_index_0_scale_req_0 : boolean;
  signal array_obj_ref_73_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_73_index_0_scale_req_1 : boolean;
  signal array_obj_ref_73_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_73_index_sum_1_req_0 : boolean;
  signal array_obj_ref_73_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_73_index_sum_1_req_1 : boolean;
  signal array_obj_ref_73_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_73_index_offset_req_0 : boolean;
  signal array_obj_ref_73_index_offset_ack_0 : boolean;
  signal array_obj_ref_73_index_offset_req_1 : boolean;
  signal array_obj_ref_73_index_offset_ack_1 : boolean;
  signal addr_of_74_final_reg_req_0 : boolean;
  signal addr_of_74_final_reg_ack_0 : boolean;
  signal addr_of_74_final_reg_req_1 : boolean;
  signal addr_of_74_final_reg_ack_1 : boolean;
  signal ptr_deref_77_store_0_req_0 : boolean;
  signal ptr_deref_77_store_0_ack_0 : boolean;
  signal ptr_deref_77_store_0_req_1 : boolean;
  signal ptr_deref_77_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeModule1_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 104) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= index;
  index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= address;
  address_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(103 downto 40) <= data;
  data_buffer <= in_buffer_data_out(103 downto 40);
  in_buffer_data_in(tag_length + 103 downto 104) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 103 downto 104);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 8,1 => 8,2 => 8,3 => 1,4 => 8);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 8);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= index_update_enable & address_update_enable & data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeModule1_CP_329_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeModule1_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= done_buffer;
  done <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule1_CP_329_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  done_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "done_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_done_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => done_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 8,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeModule1_CP_329_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule1_CP_329_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeModule1_CP_329: Block -- control-path 
    signal writeModule1_CP_329_elements: BooleanArray(36 downto 0);
    -- 
  begin -- 
    writeModule1_CP_329_elements(0) <= writeModule1_CP_329_start;
    writeModule1_CP_329_symbol <= writeModule1_CP_329_elements(36);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	15 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	27 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	18 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/$entry
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resized_0
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_computed_0
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resized_2
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scaled_2
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_computed_2
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resize_2/$entry
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resize_2/$exit
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resize_2/index_resize_req
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_resize_2/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_2/$entry
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_2/$exit
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_2/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_2/scale_rename_ack
      -- 
    writeModule1_CP_329_elements(1) <= writeModule1_CP_329_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	9 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	32 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_75_to_assign_stmt_84/index_update_enable
      -- CP-element group 2: 	 assign_stmt_75_to_assign_stmt_84/index_update_enable_out
      -- 
    writeModule1_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(29) & writeModule1_CP_329_elements(9);
      gj_writeModule1_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	16 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	33 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_75_to_assign_stmt_84/address_update_enable
      -- CP-element group 3: 	 assign_stmt_75_to_assign_stmt_84/address_update_enable_out
      -- 
    writeModule1_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_329_elements(16);
      gj_writeModule1_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	25 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	34 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_75_to_assign_stmt_84/data_update_enable
      -- CP-element group 4: 	 assign_stmt_75_to_assign_stmt_84/data_update_enable_out
      -- 
    writeModule1_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_329_elements(25);
      gj_writeModule1_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	35 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	28 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_75_to_assign_stmt_84/done_update_enable
      -- CP-element group 5: 	 assign_stmt_75_to_assign_stmt_84/done_update_enable_in
      -- 
    writeModule1_CP_329_elements(5) <= writeModule1_CP_329_elements(35);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	21 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_sample_start_
      -- CP-element group 6: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_request/$entry
      -- CP-element group 6: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_request/req
      -- 
    req_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(6), ack => addr_of_74_final_reg_req_0); -- 
    writeModule1_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(8) & writeModule1_CP_329_elements(21);
      gj_writeModule1_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	22 
    -- CP-element group 7: 	25 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	22 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_update_start_
      -- CP-element group 7: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_complete/$entry
      -- CP-element group 7: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_complete/req
      -- 
    req_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(7), ack => addr_of_74_final_reg_req_1); -- 
    writeModule1_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(1) & writeModule1_CP_329_elements(22) & writeModule1_CP_329_elements(25);
      gj_writeModule1_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	17 
    -- CP-element group 8: 	20 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_root_address_calculated
      -- CP-element group 8: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_offset_calculated
      -- CP-element group 8: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_base_plus_offset/$entry
      -- CP-element group 8: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_base_plus_offset/$exit
      -- CP-element group 8: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_base_plus_offset/sum_rename_ack
      -- 
    writeModule1_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(17) & writeModule1_CP_329_elements(20);
      gj_writeModule1_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	13 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	2 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scaled_0
      -- 
    writeModule1_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(13) & writeModule1_CP_329_elements(16);
      gj_writeModule1_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_sample_start
      -- CP-element group 10: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_Sample/rr
      -- 
    rr_364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(10), ack => array_obj_ref_73_index_0_scale_req_0); -- 
    writeModule1_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(1) & writeModule1_CP_329_elements(12);
      gj_writeModule1_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_update_start
      -- CP-element group 11: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_Update/$entry
      -- CP-element group 11: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_Update/cr
      -- 
    cr_369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(11), ack => array_obj_ref_73_index_0_scale_req_1); -- 
    writeModule1_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(1) & writeModule1_CP_329_elements(13);
      gj_writeModule1_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_sample_complete
      -- CP-element group 12: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_Sample/ra
      -- 
    ra_365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_73_index_0_scale_ack_0, ack => writeModule1_CP_329_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_update_complete
      -- CP-element group 13: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_Update/$exit
      -- CP-element group 13: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_index_scale_0_Update/ca
      -- 
    ca_370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_73_index_0_scale_ack_1, ack => writeModule1_CP_329_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_sample_start
      -- CP-element group 14: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_Sample/rr
      -- 
    rr_391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(14), ack => array_obj_ref_73_index_sum_1_req_0); -- 
    writeModule1_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 8,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(9) & writeModule1_CP_329_elements(1) & writeModule1_CP_329_elements(16);
      gj_writeModule1_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	1 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_update_start
      -- CP-element group 15: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_Update/$entry
      -- CP-element group 15: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_Update/cr
      -- 
    cr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(15), ack => array_obj_ref_73_index_sum_1_req_1); -- 
    writeModule1_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(1) & writeModule1_CP_329_elements(17) & writeModule1_CP_329_elements(19);
      gj_writeModule1_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	9 
    -- CP-element group 16: 	3 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_sample_complete
      -- CP-element group 16: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_Sample/ra
      -- 
    ra_392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_73_index_sum_1_ack_0, ack => writeModule1_CP_329_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	8 
    -- CP-element group 17: 	19 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_update_complete
      -- CP-element group 17: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_Update/$exit
      -- CP-element group 17: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_partial_sum_1_Update/ca
      -- CP-element group 17: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_Sample/$entry
      -- CP-element group 17: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_Sample/req
      -- 
    ca_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_73_index_sum_1_ack_1, ack => writeModule1_CP_329_elements(17)); -- 
    req_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(17), ack => array_obj_ref_73_index_offset_req_0); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_update_start
      -- CP-element group 18: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_Update/$entry
      -- CP-element group 18: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_Update/req
      -- 
    req_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(18), ack => array_obj_ref_73_index_offset_req_1); -- 
    writeModule1_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(1) & writeModule1_CP_329_elements(8) & writeModule1_CP_329_elements(21);
      gj_writeModule1_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	31 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_sample_complete
      -- CP-element group 19: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_Sample/ack
      -- 
    ack_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_73_index_offset_ack_0, ack => writeModule1_CP_329_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	8 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_Update/$exit
      -- CP-element group 20: 	 assign_stmt_75_to_assign_stmt_84/array_obj_ref_73_final_index_sum_regn_Update/ack
      -- 
    ack_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_73_index_offset_ack_1, ack => writeModule1_CP_329_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_sample_completed_
      -- CP-element group 21: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_request/$exit
      -- CP-element group 21: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_request/ack
      -- 
    ack_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_74_final_reg_ack_0, ack => writeModule1_CP_329_elements(21)); -- 
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	7 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	7 
    -- CP-element group 22:  members (19) 
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_update_completed_
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_complete/$exit
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/addr_of_74_complete/ack
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_address_calculated
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_word_address_calculated
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_root_address_calculated
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_address_resized
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_addr_resize/$entry
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_addr_resize/$exit
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_addr_resize/base_resize_req
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_addr_resize/base_resize_ack
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_plus_offset/$entry
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_plus_offset/$exit
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_plus_offset/sum_rename_req
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_base_plus_offset/sum_rename_ack
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_word_addrgen/$entry
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_word_addrgen/$exit
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_word_addrgen/root_register_req
      -- CP-element group 22: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_word_addrgen/root_register_ack
      -- 
    ack_424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_74_final_reg_ack_1, ack => writeModule1_CP_329_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: 	1 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_sample_start_
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/$entry
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/ptr_deref_77_Split/$entry
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/ptr_deref_77_Split/$exit
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/ptr_deref_77_Split/split_req
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/ptr_deref_77_Split/split_ack
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/word_access_start/$entry
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/word_access_start/word_0/rr
      -- 
    rr_462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(23), ack => ptr_deref_77_store_0_req_0); -- 
    writeModule1_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 8,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(22) & writeModule1_CP_329_elements(1) & writeModule1_CP_329_elements(25);
      gj_writeModule1_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_update_start_
      -- CP-element group 24: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Update/$entry
      -- CP-element group 24: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Update/word_access_complete/$entry
      -- CP-element group 24: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Update/word_access_complete/word_0/$entry
      -- CP-element group 24: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Update/word_access_complete/word_0/cr
      -- 
    cr_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(24), ack => ptr_deref_77_store_0_req_1); -- 
    writeModule1_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_329_elements(26);
      gj_writeModule1_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: 	7 
    -- CP-element group 25: 	4 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_sample_completed_
      -- CP-element group 25: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/word_access_start/$exit
      -- CP-element group 25: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Sample/word_access_start/word_0/ra
      -- 
    ra_463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_77_store_0_ack_0, ack => writeModule1_CP_329_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_update_completed_
      -- CP-element group 26: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Update/$exit
      -- CP-element group 26: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Update/word_access_complete/$exit
      -- CP-element group 26: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 assign_stmt_75_to_assign_stmt_84/ptr_deref_77_Update/word_access_complete/word_0/ca
      -- 
    ca_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_77_store_0_ack_1, ack => writeModule1_CP_329_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	1 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_sample_start_
      -- CP-element group 27: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_Sample/rr
      -- 
    rr_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(27), ack => BITSEL_u8_u1_83_inst_req_0); -- 
    writeModule1_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(1) & writeModule1_CP_329_elements(29);
      gj_writeModule1_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	5 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_update_start_
      -- CP-element group 28: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_Update/$entry
      -- CP-element group 28: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_Update/cr
      -- 
    cr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_329_elements(28), ack => BITSEL_u8_u1_83_inst_req_1); -- 
    writeModule1_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(5) & writeModule1_CP_329_elements(30);
      gj_writeModule1_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: 	2 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_sample_completed_
      -- CP-element group 29: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_Sample/$exit
      -- CP-element group 29: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_Sample/ra
      -- 
    ra_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u8_u1_83_inst_ack_0, ack => writeModule1_CP_329_elements(29)); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_update_completed_
      -- CP-element group 30: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_Update/$exit
      -- CP-element group 30: 	 assign_stmt_75_to_assign_stmt_84/BITSEL_u8_u1_83_Update/ca
      -- 
    ca_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u8_u1_83_inst_ack_1, ack => writeModule1_CP_329_elements(30)); -- 
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	12 
    -- CP-element group 31: 	19 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 assign_stmt_75_to_assign_stmt_84/$exit
      -- 
    writeModule1_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 8,1 => 8,2 => 8,3 => 8,4 => 8);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= writeModule1_CP_329_elements(16) & writeModule1_CP_329_elements(26) & writeModule1_CP_329_elements(30) & writeModule1_CP_329_elements(12) & writeModule1_CP_329_elements(19);
      gj_writeModule1_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_329_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  place  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 index_update_enable
      -- 
    writeModule1_CP_329_elements(32) <= writeModule1_CP_329_elements(2);
    -- CP-element group 33:  place  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	3 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 address_update_enable
      -- 
    writeModule1_CP_329_elements(33) <= writeModule1_CP_329_elements(3);
    -- CP-element group 34:  place  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	4 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 data_update_enable
      -- 
    writeModule1_CP_329_elements(34) <= writeModule1_CP_329_elements(4);
    -- CP-element group 35:  place  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	5 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 done_update_enable
      -- 
    -- CP-element group 36:  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	31 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 $exit
      -- 
    writeModule1_CP_329_elements(36) <= writeModule1_CP_329_elements(31);
    --  hookup: inputs to control-path 
    writeModule1_CP_329_elements(35) <= done_update_enable;
    -- hookup: output from control-path 
    index_update_enable <= writeModule1_CP_329_elements(32);
    address_update_enable <= writeModule1_CP_329_elements(33);
    data_update_enable <= writeModule1_CP_329_elements(34);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_address_72_resized : std_logic_vector(14 downto 0);
    signal R_address_72_scaled : std_logic_vector(14 downto 0);
    signal array_obj_ref_73_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_73_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_73_index_partial_sum_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_73_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_73_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_73_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_73_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_73_root_address : std_logic_vector(14 downto 0);
    signal konst_82_wire_constant : std_logic_vector(7 downto 0);
    signal ptr_75 : std_logic_vector(31 downto 0);
    signal ptr_deref_77_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_77_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_77_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_77_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_77_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_77_word_offset_0 : std_logic_vector(14 downto 0);
    signal type_cast_69_resized : std_logic_vector(14 downto 0);
    signal type_cast_69_scaled : std_logic_vector(14 downto 0);
    signal type_cast_69_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_73_constant_part_of_offset <= "000000000000000";
    array_obj_ref_73_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_73_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_73_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_73_resized_base_address <= "000000000000000";
    konst_82_wire_constant <= "00000000";
    ptr_deref_77_word_offset_0 <= "000000000000000";
    addr_of_74_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_74_final_reg_req_0;
      addr_of_74_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_74_final_reg_req_1;
      addr_of_74_final_reg_ack_1<= rack(0);
      addr_of_74_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_74_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_73_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_75,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_69_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := index_buffer(7 downto 0);
      type_cast_69_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_73_index_0_resize
    process(type_cast_69_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_69_wire;
      ov := iv(14 downto 0);
      type_cast_69_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_73_index_2_rename
    process(R_address_72_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_72_resized;
      ov(14 downto 0) := iv;
      R_address_72_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_73_index_2_resize
    process(address_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_buffer;
      ov := iv(14 downto 0);
      R_address_72_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_73_root_address_inst
    process(array_obj_ref_73_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_73_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_73_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_addr_0
    process(ptr_deref_77_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_77_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_77_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_base_resize
    process(ptr_75) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_75;
      ov := iv(14 downto 0);
      ptr_deref_77_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_gather_scatter
    process(data_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := data_buffer;
      ov(63 downto 0) := iv;
      ptr_deref_77_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_root_address_inst
    process(ptr_deref_77_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_77_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_77_root_address <= ov(14 downto 0);
      --
    end process;
    -- shared split operator group (0) : BITSEL_u8_u1_83_inst 
    ApBitsel_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= index_buffer;
      done_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= BITSEL_u8_u1_83_inst_req_0;
      BITSEL_u8_u1_83_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= BITSEL_u8_u1_83_inst_req_1;
      BITSEL_u8_u1_83_inst_ack_1 <= ackR_unguarded(0);
      ApBitsel_group_0_gI: SplitGuardInterface generic map(name => "ApBitsel_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApBitsel",
          name => "ApBitsel_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_73_index_0_scale 
    ApIntMul_group_1: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_69_resized;
      type_cast_69_scaled <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_73_index_0_scale_req_0;
      array_obj_ref_73_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_73_index_0_scale_req_1;
      array_obj_ref_73_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_1_gI: SplitGuardInterface generic map(name => "ApIntMul_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "100000000000000",
          constant_width => 15,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_73_index_offset 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= array_obj_ref_73_index_partial_sum_1;
      array_obj_ref_73_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_73_index_offset_req_0;
      array_obj_ref_73_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_73_index_offset_req_1;
      array_obj_ref_73_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "000000000000000",
          constant_width => 15,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_73_index_sum_1 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_72_scaled & type_cast_69_scaled;
      array_obj_ref_73_index_partial_sum_1 <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_73_index_sum_1_req_0;
      array_obj_ref_73_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_73_index_sum_1_req_1;
      array_obj_ref_73_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 15, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared store operator group (0) : ptr_deref_77_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(14 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 8);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_77_store_0_req_0;
      ptr_deref_77_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_77_store_0_req_1;
      ptr_deref_77_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_77_word_address_0;
      data_in <= ptr_deref_77_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 15,
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(14 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end writeModule1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(14 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(14 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    Zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    Zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    zeropad_same_call_reqs : out  std_logic_vector(0 downto 0);
    zeropad_same_call_acks : in   std_logic_vector(0 downto 0);
    zeropad_same_call_data : out  std_logic_vector(111 downto 0);
    zeropad_same_call_tag  :  out  std_logic_vector(0 downto 0);
    zeropad_same_return_reqs : out  std_logic_vector(0 downto 0);
    zeropad_same_return_acks : in   std_logic_vector(0 downto 0);
    zeropad_same_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad;
architecture zeropad_arch of zeropad is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad_CP_920_start: Boolean;
  signal zeropad_CP_920_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component zeropad_same is -- 
    generic (tag_length : integer); 
    port ( -- 
      inp_d0 : in  std_logic_vector(15 downto 0);
      inp_d1 : in  std_logic_vector(15 downto 0);
      inp_d2 : in  std_logic_vector(15 downto 0);
      out_d0 : in  std_logic_vector(15 downto 0);
      out_d1 : in  std_logic_vector(15 downto 0);
      out_d2 : in  std_logic_vector(15 downto 0);
      index1 : in  std_logic_vector(7 downto 0);
      index2 : in  std_logic_vector(7 downto 0);
      readModule1_call_reqs : out  std_logic_vector(0 downto 0);
      readModule1_call_acks : in   std_logic_vector(0 downto 0);
      readModule1_call_data : out  std_logic_vector(39 downto 0);
      readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      readModule1_return_reqs : out  std_logic_vector(0 downto 0);
      readModule1_return_acks : in   std_logic_vector(0 downto 0);
      readModule1_return_data : in   std_logic_vector(63 downto 0);
      readModule1_return_tag :  in   std_logic_vector(0 downto 0);
      writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_call_acks : in   std_logic_vector(0 downto 0);
      writeModule1_call_data : out  std_logic_vector(103 downto 0);
      writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_return_acks : in   std_logic_vector(0 downto 0);
      writeModule1_return_data : in   std_logic_vector(0 downto 0);
      writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_435_inst_ack_0 : boolean;
  signal type_cast_491_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_456_inst_ack_0 : boolean;
  signal addr_of_812_final_reg_ack_1 : boolean;
  signal type_cast_397_inst_ack_0 : boolean;
  signal if_stmt_830_branch_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_393_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_368_inst_ack_0 : boolean;
  signal type_cast_491_inst_req_1 : boolean;
  signal type_cast_945_inst_req_1 : boolean;
  signal type_cast_469_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_356_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_456_inst_req_0 : boolean;
  signal type_cast_422_inst_req_1 : boolean;
  signal type_cast_422_inst_ack_1 : boolean;
  signal type_cast_915_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_418_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_356_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_418_inst_ack_0 : boolean;
  signal type_cast_435_inst_req_0 : boolean;
  signal type_cast_915_inst_req_1 : boolean;
  signal type_cast_397_inst_req_0 : boolean;
  signal type_cast_435_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_356_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_393_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_381_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_443_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_381_inst_req_0 : boolean;
  signal type_cast_372_inst_ack_1 : boolean;
  signal type_cast_372_inst_req_1 : boolean;
  signal type_cast_422_inst_req_0 : boolean;
  signal type_cast_447_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_393_inst_req_1 : boolean;
  signal type_cast_397_inst_req_1 : boolean;
  signal type_cast_447_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_431_inst_req_0 : boolean;
  signal type_cast_397_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_950_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_356_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_393_inst_ack_0 : boolean;
  signal if_stmt_830_branch_req_0 : boolean;
  signal type_cast_477_inst_req_0 : boolean;
  signal call_stmt_862_call_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_443_inst_ack_1 : boolean;
  signal type_cast_477_inst_ack_0 : boolean;
  signal type_cast_469_inst_ack_0 : boolean;
  signal call_stmt_862_call_req_1 : boolean;
  signal type_cast_447_inst_ack_0 : boolean;
  signal type_cast_360_inst_req_1 : boolean;
  signal type_cast_915_inst_ack_1 : boolean;
  signal call_stmt_862_call_req_0 : boolean;
  signal type_cast_945_inst_ack_1 : boolean;
  signal type_cast_491_inst_ack_1 : boolean;
  signal type_cast_435_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_431_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_431_inst_ack_0 : boolean;
  signal type_cast_410_inst_ack_0 : boolean;
  signal ptr_deref_815_store_0_ack_1 : boolean;
  signal type_cast_469_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_418_inst_req_0 : boolean;
  signal type_cast_360_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_368_inst_req_0 : boolean;
  signal type_cast_385_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_443_inst_req_1 : boolean;
  signal type_cast_385_inst_req_1 : boolean;
  signal type_cast_473_inst_req_1 : boolean;
  signal type_cast_469_inst_req_1 : boolean;
  signal type_cast_473_inst_ack_1 : boolean;
  signal type_cast_360_inst_ack_0 : boolean;
  signal type_cast_460_inst_req_0 : boolean;
  signal type_cast_895_inst_req_0 : boolean;
  signal type_cast_385_inst_req_0 : boolean;
  signal type_cast_385_inst_ack_0 : boolean;
  signal addr_of_812_final_reg_req_1 : boolean;
  signal type_cast_473_inst_ack_0 : boolean;
  signal type_cast_422_inst_ack_0 : boolean;
  signal type_cast_473_inst_req_0 : boolean;
  signal type_cast_491_inst_req_0 : boolean;
  signal type_cast_477_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_431_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_381_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_381_inst_ack_0 : boolean;
  signal type_cast_477_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_418_inst_ack_1 : boolean;
  signal type_cast_410_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_443_inst_ack_0 : boolean;
  signal type_cast_410_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_456_inst_req_1 : boolean;
  signal type_cast_410_inst_req_0 : boolean;
  signal type_cast_460_inst_ack_1 : boolean;
  signal call_stmt_862_call_ack_0 : boolean;
  signal type_cast_372_inst_ack_0 : boolean;
  signal type_cast_372_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_406_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_406_inst_req_1 : boolean;
  signal type_cast_447_inst_req_1 : boolean;
  signal type_cast_460_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_406_inst_ack_0 : boolean;
  signal type_cast_460_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_406_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_456_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_368_inst_ack_1 : boolean;
  signal if_stmt_830_branch_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_368_inst_req_1 : boolean;
  signal type_cast_925_inst_req_0 : boolean;
  signal type_cast_360_inst_ack_1 : boolean;
  signal type_cast_925_inst_ack_0 : boolean;
  signal type_cast_895_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_962_inst_ack_0 : boolean;
  signal type_cast_866_inst_req_0 : boolean;
  signal type_cast_925_inst_req_1 : boolean;
  signal type_cast_866_inst_ack_0 : boolean;
  signal type_cast_925_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_959_inst_ack_1 : boolean;
  signal type_cast_866_inst_req_1 : boolean;
  signal type_cast_866_inst_ack_1 : boolean;
  signal type_cast_875_inst_req_0 : boolean;
  signal type_cast_875_inst_ack_0 : boolean;
  signal type_cast_935_inst_req_0 : boolean;
  signal type_cast_935_inst_ack_0 : boolean;
  signal type_cast_875_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_947_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_953_inst_req_0 : boolean;
  signal call_stmt_841_call_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_965_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_959_inst_req_0 : boolean;
  signal type_cast_875_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_959_inst_ack_0 : boolean;
  signal call_stmt_841_call_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_953_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_947_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_965_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_962_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_962_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_962_inst_req_0 : boolean;
  signal call_stmt_841_call_req_1 : boolean;
  signal call_stmt_841_call_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_968_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_965_inst_req_1 : boolean;
  signal type_cast_846_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_968_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_965_inst_ack_1 : boolean;
  signal phi_stmt_797_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_318_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_318_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_318_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_318_inst_ack_1 : boolean;
  signal type_cast_322_inst_req_0 : boolean;
  signal type_cast_322_inst_ack_0 : boolean;
  signal type_cast_322_inst_req_1 : boolean;
  signal type_cast_322_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_331_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_331_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_331_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_331_inst_ack_1 : boolean;
  signal type_cast_335_inst_req_0 : boolean;
  signal type_cast_335_inst_ack_0 : boolean;
  signal type_cast_335_inst_req_1 : boolean;
  signal type_cast_335_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_343_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_343_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_343_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_343_inst_ack_1 : boolean;
  signal type_cast_347_inst_req_0 : boolean;
  signal type_cast_347_inst_ack_0 : boolean;
  signal type_cast_347_inst_req_1 : boolean;
  signal type_cast_347_inst_ack_1 : boolean;
  signal ptr_deref_815_store_0_req_1 : boolean;
  signal type_cast_945_inst_ack_0 : boolean;
  signal type_cast_915_inst_req_0 : boolean;
  signal type_cast_495_inst_req_0 : boolean;
  signal type_cast_495_inst_ack_0 : boolean;
  signal type_cast_495_inst_req_1 : boolean;
  signal type_cast_495_inst_ack_1 : boolean;
  signal type_cast_945_inst_req_0 : boolean;
  signal call_stmt_859_call_ack_1 : boolean;
  signal type_cast_499_inst_req_0 : boolean;
  signal type_cast_499_inst_ack_0 : boolean;
  signal addr_of_812_final_reg_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_956_inst_ack_1 : boolean;
  signal type_cast_499_inst_req_1 : boolean;
  signal type_cast_499_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_950_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_950_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_950_inst_req_0 : boolean;
  signal call_stmt_859_call_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_956_inst_req_1 : boolean;
  signal if_stmt_517_branch_req_0 : boolean;
  signal if_stmt_517_branch_ack_1 : boolean;
  signal addr_of_812_final_reg_req_0 : boolean;
  signal if_stmt_517_branch_ack_0 : boolean;
  signal type_cast_885_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_959_inst_req_1 : boolean;
  signal type_cast_885_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_956_inst_ack_0 : boolean;
  signal if_stmt_532_branch_req_0 : boolean;
  signal if_stmt_532_branch_ack_1 : boolean;
  signal if_stmt_532_branch_ack_0 : boolean;
  signal type_cast_885_inst_ack_0 : boolean;
  signal type_cast_905_inst_ack_1 : boolean;
  signal call_stmt_859_call_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_956_inst_req_0 : boolean;
  signal type_cast_541_inst_req_0 : boolean;
  signal type_cast_905_inst_req_1 : boolean;
  signal type_cast_541_inst_ack_0 : boolean;
  signal type_cast_885_inst_req_0 : boolean;
  signal type_cast_541_inst_req_1 : boolean;
  signal type_cast_541_inst_ack_1 : boolean;
  signal ptr_deref_815_store_0_ack_0 : boolean;
  signal ptr_deref_815_store_0_req_0 : boolean;
  signal call_stmt_859_call_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_947_inst_ack_0 : boolean;
  signal type_cast_545_inst_req_0 : boolean;
  signal type_cast_545_inst_ack_0 : boolean;
  signal type_cast_545_inst_req_1 : boolean;
  signal type_cast_905_inst_ack_0 : boolean;
  signal type_cast_545_inst_ack_1 : boolean;
  signal type_cast_935_inst_ack_1 : boolean;
  signal type_cast_554_inst_req_0 : boolean;
  signal type_cast_905_inst_req_0 : boolean;
  signal type_cast_554_inst_ack_0 : boolean;
  signal type_cast_554_inst_req_1 : boolean;
  signal type_cast_554_inst_ack_1 : boolean;
  signal type_cast_935_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_947_inst_req_0 : boolean;
  signal type_cast_846_inst_ack_1 : boolean;
  signal type_cast_846_inst_req_1 : boolean;
  signal array_obj_ref_596_index_offset_req_0 : boolean;
  signal array_obj_ref_596_index_offset_ack_0 : boolean;
  signal array_obj_ref_596_index_offset_req_1 : boolean;
  signal array_obj_ref_596_index_offset_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_953_inst_req_1 : boolean;
  signal type_cast_846_inst_ack_0 : boolean;
  signal addr_of_597_final_reg_req_0 : boolean;
  signal type_cast_895_inst_ack_1 : boolean;
  signal addr_of_597_final_reg_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_953_inst_ack_1 : boolean;
  signal addr_of_597_final_reg_req_1 : boolean;
  signal type_cast_895_inst_req_1 : boolean;
  signal addr_of_597_final_reg_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_600_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_600_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_600_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_600_inst_ack_1 : boolean;
  signal type_cast_604_inst_req_0 : boolean;
  signal type_cast_604_inst_ack_0 : boolean;
  signal type_cast_604_inst_req_1 : boolean;
  signal type_cast_604_inst_ack_1 : boolean;
  signal phi_stmt_582_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_613_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_613_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_613_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_613_inst_ack_1 : boolean;
  signal type_cast_1028_inst_req_0 : boolean;
  signal type_cast_1028_inst_ack_0 : boolean;
  signal type_cast_617_inst_req_0 : boolean;
  signal type_cast_617_inst_ack_0 : boolean;
  signal type_cast_617_inst_req_1 : boolean;
  signal type_cast_617_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_631_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_631_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_631_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_631_inst_ack_1 : boolean;
  signal type_cast_1028_inst_req_1 : boolean;
  signal type_cast_1028_inst_ack_1 : boolean;
  signal type_cast_635_inst_req_0 : boolean;
  signal type_cast_635_inst_ack_0 : boolean;
  signal type_cast_635_inst_req_1 : boolean;
  signal type_cast_635_inst_ack_1 : boolean;
  signal phi_stmt_1022_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_649_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_649_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_649_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_649_inst_ack_1 : boolean;
  signal type_cast_653_inst_req_0 : boolean;
  signal type_cast_653_inst_ack_0 : boolean;
  signal type_cast_653_inst_req_1 : boolean;
  signal type_cast_653_inst_ack_1 : boolean;
  signal phi_stmt_1022_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_667_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_667_inst_ack_0 : boolean;
  signal type_cast_803_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_667_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_667_inst_ack_1 : boolean;
  signal type_cast_803_inst_ack_0 : boolean;
  signal type_cast_671_inst_req_0 : boolean;
  signal type_cast_671_inst_ack_0 : boolean;
  signal type_cast_671_inst_req_1 : boolean;
  signal type_cast_671_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_685_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_685_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_685_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_685_inst_ack_1 : boolean;
  signal type_cast_803_inst_req_1 : boolean;
  signal type_cast_689_inst_req_0 : boolean;
  signal type_cast_689_inst_ack_0 : boolean;
  signal type_cast_689_inst_req_1 : boolean;
  signal type_cast_689_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_703_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_703_inst_ack_0 : boolean;
  signal type_cast_803_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_703_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_703_inst_ack_1 : boolean;
  signal type_cast_707_inst_req_0 : boolean;
  signal type_cast_707_inst_ack_0 : boolean;
  signal type_cast_707_inst_req_1 : boolean;
  signal phi_stmt_797_req_1 : boolean;
  signal type_cast_707_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_721_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_721_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_721_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_721_inst_ack_1 : boolean;
  signal type_cast_725_inst_req_0 : boolean;
  signal type_cast_725_inst_ack_0 : boolean;
  signal type_cast_725_inst_req_1 : boolean;
  signal type_cast_725_inst_ack_1 : boolean;
  signal ptr_deref_733_store_0_req_0 : boolean;
  signal ptr_deref_733_store_0_ack_0 : boolean;
  signal ptr_deref_733_store_0_req_1 : boolean;
  signal ptr_deref_733_store_0_ack_1 : boolean;
  signal if_stmt_747_branch_req_0 : boolean;
  signal if_stmt_747_branch_ack_1 : boolean;
  signal if_stmt_747_branch_ack_0 : boolean;
  signal type_cast_756_inst_req_0 : boolean;
  signal type_cast_756_inst_ack_0 : boolean;
  signal type_cast_756_inst_req_1 : boolean;
  signal type_cast_756_inst_ack_1 : boolean;
  signal type_cast_760_inst_req_0 : boolean;
  signal type_cast_760_inst_ack_0 : boolean;
  signal type_cast_760_inst_req_1 : boolean;
  signal type_cast_760_inst_ack_1 : boolean;
  signal type_cast_769_inst_req_0 : boolean;
  signal type_cast_769_inst_ack_0 : boolean;
  signal type_cast_769_inst_req_1 : boolean;
  signal type_cast_769_inst_ack_1 : boolean;
  signal array_obj_ref_811_index_offset_req_0 : boolean;
  signal array_obj_ref_811_index_offset_ack_0 : boolean;
  signal array_obj_ref_811_index_offset_req_1 : boolean;
  signal array_obj_ref_811_index_offset_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_968_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_968_inst_ack_1 : boolean;
  signal phi_stmt_582_ack_0 : boolean;
  signal phi_stmt_582_req_1 : boolean;
  signal type_cast_588_inst_ack_1 : boolean;
  signal type_cast_588_inst_req_1 : boolean;
  signal type_cast_588_inst_ack_0 : boolean;
  signal type_cast_588_inst_req_0 : boolean;
  signal phi_stmt_1022_req_0 : boolean;
  signal if_stmt_972_branch_req_0 : boolean;
  signal if_stmt_972_branch_ack_1 : boolean;
  signal if_stmt_972_branch_ack_0 : boolean;
  signal type_cast_981_inst_req_0 : boolean;
  signal type_cast_981_inst_ack_0 : boolean;
  signal type_cast_981_inst_req_1 : boolean;
  signal type_cast_981_inst_ack_1 : boolean;
  signal type_cast_985_inst_req_0 : boolean;
  signal type_cast_985_inst_ack_0 : boolean;
  signal type_cast_985_inst_req_1 : boolean;
  signal type_cast_985_inst_ack_1 : boolean;
  signal type_cast_994_inst_req_0 : boolean;
  signal type_cast_994_inst_ack_0 : boolean;
  signal type_cast_994_inst_req_1 : boolean;
  signal type_cast_994_inst_ack_1 : boolean;
  signal array_obj_ref_1036_index_offset_req_0 : boolean;
  signal array_obj_ref_1036_index_offset_ack_0 : boolean;
  signal array_obj_ref_1036_index_offset_req_1 : boolean;
  signal array_obj_ref_1036_index_offset_ack_1 : boolean;
  signal addr_of_1037_final_reg_req_0 : boolean;
  signal addr_of_1037_final_reg_ack_0 : boolean;
  signal addr_of_1037_final_reg_req_1 : boolean;
  signal addr_of_1037_final_reg_ack_1 : boolean;
  signal phi_stmt_797_ack_0 : boolean;
  signal ptr_deref_1041_load_0_req_0 : boolean;
  signal ptr_deref_1041_load_0_ack_0 : boolean;
  signal ptr_deref_1041_load_0_req_1 : boolean;
  signal ptr_deref_1041_load_0_ack_1 : boolean;
  signal type_cast_1045_inst_req_0 : boolean;
  signal type_cast_1045_inst_ack_0 : boolean;
  signal type_cast_1045_inst_req_1 : boolean;
  signal type_cast_1045_inst_ack_1 : boolean;
  signal type_cast_1055_inst_req_0 : boolean;
  signal type_cast_1055_inst_ack_0 : boolean;
  signal type_cast_1055_inst_req_1 : boolean;
  signal type_cast_1055_inst_ack_1 : boolean;
  signal type_cast_1065_inst_req_0 : boolean;
  signal type_cast_1065_inst_ack_0 : boolean;
  signal type_cast_1065_inst_req_1 : boolean;
  signal type_cast_1065_inst_ack_1 : boolean;
  signal type_cast_1075_inst_req_0 : boolean;
  signal type_cast_1075_inst_ack_0 : boolean;
  signal type_cast_1075_inst_req_1 : boolean;
  signal type_cast_1075_inst_ack_1 : boolean;
  signal type_cast_1085_inst_req_0 : boolean;
  signal type_cast_1085_inst_ack_0 : boolean;
  signal type_cast_1085_inst_req_1 : boolean;
  signal type_cast_1085_inst_ack_1 : boolean;
  signal type_cast_1095_inst_req_0 : boolean;
  signal type_cast_1095_inst_ack_0 : boolean;
  signal type_cast_1095_inst_req_1 : boolean;
  signal type_cast_1095_inst_ack_1 : boolean;
  signal type_cast_1105_inst_req_0 : boolean;
  signal type_cast_1105_inst_ack_0 : boolean;
  signal type_cast_1105_inst_req_1 : boolean;
  signal type_cast_1105_inst_ack_1 : boolean;
  signal type_cast_1115_inst_req_0 : boolean;
  signal type_cast_1115_inst_ack_0 : boolean;
  signal type_cast_1115_inst_req_1 : boolean;
  signal type_cast_1115_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1117_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1117_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1117_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1117_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1120_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1120_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1120_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1120_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1123_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1123_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1123_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1123_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1126_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1126_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1126_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1126_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1129_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1129_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1129_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1129_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1132_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1132_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1132_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1132_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1135_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1135_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1135_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1135_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1138_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1138_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1138_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1138_inst_ack_1 : boolean;
  signal if_stmt_1152_branch_req_0 : boolean;
  signal if_stmt_1152_branch_ack_1 : boolean;
  signal if_stmt_1152_branch_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad_CP_920_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad_CP_920_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad_CP_920_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad_CP_920_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad_CP_920: Block -- control-path 
    signal zeropad_CP_920_elements: BooleanArray(263 downto 0);
    -- 
  begin -- 
    zeropad_CP_920_elements(0) <= zeropad_CP_920_start;
    zeropad_CP_920_symbol <= zeropad_CP_920_elements(263);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	54 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	66 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	51 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	63 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0:  members (62) 
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_316/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/branch_block_stmt_316__entry__
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516__entry__
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_update_start_
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_Update/cr
      -- 
    cr_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_491_inst_req_1); -- 
    cr_1241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_422_inst_req_1); -- 
    cr_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_372_inst_req_1); -- 
    cr_1185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_397_inst_req_1); -- 
    cr_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_360_inst_req_1); -- 
    cr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_435_inst_req_1); -- 
    cr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_385_inst_req_1); -- 
    cr_1353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_473_inst_req_1); -- 
    cr_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_469_inst_req_1); -- 
    cr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_477_inst_req_1); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_410_inst_req_1); -- 
    cr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_447_inst_req_1); -- 
    cr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_460_inst_req_1); -- 
    rr_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => RPIPE_Zeropad_input_pipe_318_inst_req_0); -- 
    cr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_322_inst_req_1); -- 
    cr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_335_inst_req_1); -- 
    cr_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_347_inst_req_1); -- 
    cr_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_495_inst_req_1); -- 
    cr_1409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(0), ack => type_cast_499_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_update_start_
      -- CP-element group 1: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_Update/cr
      -- 
    ra_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_318_inst_ack_0, ack => zeropad_CP_920_elements(1)); -- 
    cr_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(1), ack => RPIPE_Zeropad_input_pipe_318_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_318_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_Sample/rr
      -- 
    ca_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_318_inst_ack_1, ack => zeropad_CP_920_elements(2)); -- 
    rr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(2), ack => type_cast_322_inst_req_0); -- 
    rr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(2), ack => RPIPE_Zeropad_input_pipe_331_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_Sample/ra
      -- 
    ra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_0, ack => zeropad_CP_920_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	49 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_322_Update/ca
      -- 
    ca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_1, ack => zeropad_CP_920_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_update_start_
      -- CP-element group 5: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_Update/cr
      -- 
    ra_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_331_inst_ack_0, ack => zeropad_CP_920_elements(5)); -- 
    cr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(5), ack => RPIPE_Zeropad_input_pipe_331_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_331_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_Sample/rr
      -- 
    ca_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_331_inst_ack_1, ack => zeropad_CP_920_elements(6)); -- 
    rr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(6), ack => type_cast_335_inst_req_0); -- 
    rr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(6), ack => RPIPE_Zeropad_input_pipe_343_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_Sample/ra
      -- 
    ra_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_335_inst_ack_0, ack => zeropad_CP_920_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	49 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_335_Update/ca
      -- 
    ca_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_335_inst_ack_1, ack => zeropad_CP_920_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_update_start_
      -- CP-element group 9: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_Update/cr
      -- 
    ra_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_343_inst_ack_0, ack => zeropad_CP_920_elements(9)); -- 
    cr_1059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(9), ack => RPIPE_Zeropad_input_pipe_343_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_343_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_Sample/rr
      -- 
    ca_1060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_343_inst_ack_1, ack => zeropad_CP_920_elements(10)); -- 
    rr_1082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(10), ack => RPIPE_Zeropad_input_pipe_356_inst_req_0); -- 
    rr_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(10), ack => type_cast_347_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_Sample/ra
      -- 
    ra_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_347_inst_ack_0, ack => zeropad_CP_920_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	52 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_347_Update/ca
      -- 
    ca_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_347_inst_ack_1, ack => zeropad_CP_920_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_update_start_
      -- CP-element group 13: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_sample_completed_
      -- 
    ra_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_356_inst_ack_0, ack => zeropad_CP_920_elements(13)); -- 
    cr_1087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(13), ack => RPIPE_Zeropad_input_pipe_356_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_356_update_completed_
      -- 
    ca_1088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_356_inst_ack_1, ack => zeropad_CP_920_elements(14)); -- 
    rr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(14), ack => RPIPE_Zeropad_input_pipe_368_inst_req_0); -- 
    rr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(14), ack => type_cast_360_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_Sample/ra
      -- 
    ra_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_0, ack => zeropad_CP_920_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	52 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_360_Update/ca
      -- 
    ca_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_1, ack => zeropad_CP_920_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_update_start_
      -- CP-element group 17: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_Update/cr
      -- 
    ra_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_368_inst_ack_0, ack => zeropad_CP_920_elements(17)); -- 
    cr_1115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(17), ack => RPIPE_Zeropad_input_pipe_368_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_368_Update/ca
      -- 
    ca_1116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_368_inst_ack_1, ack => zeropad_CP_920_elements(18)); -- 
    rr_1124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(18), ack => type_cast_372_inst_req_0); -- 
    rr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(18), ack => RPIPE_Zeropad_input_pipe_381_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_sample_completed_
      -- 
    ra_1125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_372_inst_ack_0, ack => zeropad_CP_920_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	55 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_372_update_completed_
      -- 
    ca_1130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_372_inst_ack_1, ack => zeropad_CP_920_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_update_start_
      -- CP-element group 21: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_Sample/$exit
      -- 
    ra_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_381_inst_ack_0, ack => zeropad_CP_920_elements(21)); -- 
    cr_1143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(21), ack => RPIPE_Zeropad_input_pipe_381_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_381_update_completed_
      -- 
    ca_1144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_381_inst_ack_1, ack => zeropad_CP_920_elements(22)); -- 
    rr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(22), ack => type_cast_385_inst_req_0); -- 
    rr_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(22), ack => RPIPE_Zeropad_input_pipe_393_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_Sample/ra
      -- 
    ra_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_385_inst_ack_0, ack => zeropad_CP_920_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	55 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_385_update_completed_
      -- 
    ca_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_385_inst_ack_1, ack => zeropad_CP_920_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_update_start_
      -- CP-element group 25: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_Update/$entry
      -- 
    ra_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_393_inst_ack_0, ack => zeropad_CP_920_elements(25)); -- 
    cr_1171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(25), ack => RPIPE_Zeropad_input_pipe_393_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_393_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_Sample/$entry
      -- 
    ca_1172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_393_inst_ack_1, ack => zeropad_CP_920_elements(26)); -- 
    rr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(26), ack => type_cast_397_inst_req_0); -- 
    rr_1194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(26), ack => RPIPE_Zeropad_input_pipe_406_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_sample_completed_
      -- 
    ra_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_397_inst_ack_0, ack => zeropad_CP_920_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	58 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_397_update_completed_
      -- 
    ca_1186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_397_inst_ack_1, ack => zeropad_CP_920_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_update_start_
      -- CP-element group 29: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_Sample/$exit
      -- 
    ra_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_406_inst_ack_0, ack => zeropad_CP_920_elements(29)); -- 
    cr_1199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(29), ack => RPIPE_Zeropad_input_pipe_406_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_406_Update/$exit
      -- 
    ca_1200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_406_inst_ack_1, ack => zeropad_CP_920_elements(30)); -- 
    rr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(30), ack => type_cast_410_inst_req_0); -- 
    rr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(30), ack => RPIPE_Zeropad_input_pipe_418_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_sample_completed_
      -- 
    ra_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_410_inst_ack_0, ack => zeropad_CP_920_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	58 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_410_update_completed_
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_410_inst_ack_1, ack => zeropad_CP_920_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_update_start_
      -- CP-element group 33: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_Update/$entry
      -- 
    ra_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_418_inst_ack_0, ack => zeropad_CP_920_elements(33)); -- 
    cr_1227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(33), ack => RPIPE_Zeropad_input_pipe_418_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_418_Update/ca
      -- 
    ca_1228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_418_inst_ack_1, ack => zeropad_CP_920_elements(34)); -- 
    rr_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(34), ack => type_cast_422_inst_req_0); -- 
    rr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(34), ack => RPIPE_Zeropad_input_pipe_431_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_Sample/ra
      -- 
    ra_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_422_inst_ack_0, ack => zeropad_CP_920_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	61 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_422_Update/$exit
      -- 
    ca_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_422_inst_ack_1, ack => zeropad_CP_920_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_update_start_
      -- CP-element group 37: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_Update/cr
      -- 
    ra_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_431_inst_ack_0, ack => zeropad_CP_920_elements(37)); -- 
    cr_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(37), ack => RPIPE_Zeropad_input_pipe_431_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_431_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_sample_start_
      -- 
    ca_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_431_inst_ack_1, ack => zeropad_CP_920_elements(38)); -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(38), ack => type_cast_435_inst_req_0); -- 
    rr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(38), ack => RPIPE_Zeropad_input_pipe_443_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_sample_completed_
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_435_inst_ack_0, ack => zeropad_CP_920_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	61 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_435_update_completed_
      -- 
    ca_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_435_inst_ack_1, ack => zeropad_CP_920_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_update_start_
      -- CP-element group 41: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_Sample/ra
      -- 
    ra_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_443_inst_ack_0, ack => zeropad_CP_920_elements(41)); -- 
    cr_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(41), ack => RPIPE_Zeropad_input_pipe_443_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_443_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_Sample/$entry
      -- 
    ca_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_443_inst_ack_1, ack => zeropad_CP_920_elements(42)); -- 
    rr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(42), ack => type_cast_447_inst_req_0); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(42), ack => RPIPE_Zeropad_input_pipe_456_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_sample_completed_
      -- 
    ra_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_447_inst_ack_0, ack => zeropad_CP_920_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	64 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_447_Update/$exit
      -- 
    ca_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_447_inst_ack_1, ack => zeropad_CP_920_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_update_start_
      -- CP-element group 45: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_Update/cr
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_456_inst_ack_0, ack => zeropad_CP_920_elements(45)); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(45), ack => RPIPE_Zeropad_input_pipe_456_inst_req_1); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/RPIPE_Zeropad_input_pipe_456_Update/ca
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_456_inst_ack_1, ack => zeropad_CP_920_elements(46)); -- 
    rr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(46), ack => type_cast_460_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_Sample/ra
      -- 
    ra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_460_inst_ack_0, ack => zeropad_CP_920_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	64 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_460_Update/$exit
      -- 
    ca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_460_inst_ack_1, ack => zeropad_CP_920_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	4 
    -- CP-element group 49: 	8 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_sample_start_
      -- 
    rr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(49), ack => type_cast_469_inst_req_0); -- 
    zeropad_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(4) & zeropad_CP_920_elements(8);
      gj_zeropad_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_Sample/ra
      -- 
    ra_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_469_inst_ack_0, ack => zeropad_CP_920_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	0 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	67 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_469_Update/ca
      -- 
    ca_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_469_inst_ack_1, ack => zeropad_CP_920_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	16 
    -- CP-element group 52: 	12 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_sample_start_
      -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(52), ack => type_cast_473_inst_req_0); -- 
    zeropad_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(16) & zeropad_CP_920_elements(12);
      gj_zeropad_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_sample_completed_
      -- 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_0, ack => zeropad_CP_920_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	67 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_473_update_completed_
      -- 
    ca_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_1, ack => zeropad_CP_920_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	20 
    -- CP-element group 55: 	24 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_sample_start_
      -- 
    rr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(55), ack => type_cast_477_inst_req_0); -- 
    zeropad_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(20) & zeropad_CP_920_elements(24);
      gj_zeropad_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_sample_completed_
      -- 
    ra_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_477_inst_ack_0, ack => zeropad_CP_920_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	67 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_477_Update/ca
      -- 
    ca_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_477_inst_ack_1, ack => zeropad_CP_920_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	28 
    -- CP-element group 58: 	32 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_sample_start_
      -- 
    rr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(58), ack => type_cast_491_inst_req_0); -- 
    zeropad_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(28) & zeropad_CP_920_elements(32);
      gj_zeropad_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_Sample/ra
      -- CP-element group 59: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_Sample/$exit
      -- 
    ra_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_491_inst_ack_0, ack => zeropad_CP_920_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	67 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_491_Update/ca
      -- 
    ca_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_491_inst_ack_1, ack => zeropad_CP_920_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	36 
    -- CP-element group 61: 	40 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_Sample/rr
      -- 
    rr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(61), ack => type_cast_495_inst_req_0); -- 
    zeropad_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(36) & zeropad_CP_920_elements(40);
      gj_zeropad_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_Sample/ra
      -- 
    ra_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_495_inst_ack_0, ack => zeropad_CP_920_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	0 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	67 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_495_Update/ca
      -- 
    ca_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_495_inst_ack_1, ack => zeropad_CP_920_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	44 
    -- CP-element group 64: 	48 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_Sample/rr
      -- 
    rr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(64), ack => type_cast_499_inst_req_0); -- 
    zeropad_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(44) & zeropad_CP_920_elements(48);
      gj_zeropad_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_Sample/ra
      -- 
    ra_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_499_inst_ack_0, ack => zeropad_CP_920_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	0 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/type_cast_499_Update/ca
      -- 
    ca_1410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_499_inst_ack_1, ack => zeropad_CP_920_elements(66)); -- 
    -- CP-element group 67:  branch  join  transition  place  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	54 
    -- CP-element group 67: 	66 
    -- CP-element group 67: 	51 
    -- CP-element group 67: 	60 
    -- CP-element group 67: 	63 
    -- CP-element group 67: 	57 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (10) 
      -- CP-element group 67: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516__exit__
      -- CP-element group 67: 	 branch_block_stmt_316/if_stmt_517__entry__
      -- CP-element group 67: 	 branch_block_stmt_316/assign_stmt_319_to_assign_stmt_516/$exit
      -- CP-element group 67: 	 branch_block_stmt_316/if_stmt_517_dead_link/$entry
      -- CP-element group 67: 	 branch_block_stmt_316/if_stmt_517_eval_test/$entry
      -- CP-element group 67: 	 branch_block_stmt_316/if_stmt_517_eval_test/$exit
      -- CP-element group 67: 	 branch_block_stmt_316/if_stmt_517_eval_test/branch_req
      -- CP-element group 67: 	 branch_block_stmt_316/R_cmp296_518_place
      -- CP-element group 67: 	 branch_block_stmt_316/if_stmt_517_if_link/$entry
      -- CP-element group 67: 	 branch_block_stmt_316/if_stmt_517_else_link/$entry
      -- 
    branch_req_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(67), ack => if_stmt_517_branch_req_0); -- 
    zeropad_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(54) & zeropad_CP_920_elements(66) & zeropad_CP_920_elements(51) & zeropad_CP_920_elements(60) & zeropad_CP_920_elements(63) & zeropad_CP_920_elements(57);
      gj_zeropad_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	72 
    -- CP-element group 68: 	73 
    -- CP-element group 68: 	74 
    -- CP-element group 68: 	75 
    -- CP-element group 68: 	76 
    -- CP-element group 68: 	77 
    -- CP-element group 68:  members (30) 
      -- CP-element group 68: 	 branch_block_stmt_316/merge_stmt_538__exit__
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579__entry__
      -- CP-element group 68: 	 branch_block_stmt_316/if_stmt_517_if_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_316/if_stmt_517_if_link/if_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_316/entry_bbx_xnph298
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_update_start_
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_update_start_
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_update_start_
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_316/merge_stmt_538_PhiAck/dummy
      -- CP-element group 68: 	 branch_block_stmt_316/merge_stmt_538_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_316/merge_stmt_538_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/entry_bbx_xnph298_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_316/entry_bbx_xnph298_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_316/merge_stmt_538_PhiReqMerge
      -- 
    if_choice_transition_1423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_517_branch_ack_1, ack => zeropad_CP_920_elements(68)); -- 
    rr_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(68), ack => type_cast_541_inst_req_0); -- 
    cr_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(68), ack => type_cast_541_inst_req_1); -- 
    rr_1476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(68), ack => type_cast_545_inst_req_0); -- 
    cr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(68), ack => type_cast_545_inst_req_1); -- 
    rr_1490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(68), ack => type_cast_554_inst_req_0); -- 
    cr_1495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(68), ack => type_cast_554_inst_req_1); -- 
    -- CP-element group 69:  transition  place  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	243 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_316/if_stmt_517_else_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_316/if_stmt_517_else_link/else_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_316/entry_forx_xcond119x_xpreheader
      -- CP-element group 69: 	 branch_block_stmt_316/entry_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_316/entry_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_1427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_517_branch_ack_0, ack => zeropad_CP_920_elements(69)); -- 
    -- CP-element group 70:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	243 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	125 
    -- CP-element group 70: 	126 
    -- CP-element group 70: 	121 
    -- CP-element group 70: 	122 
    -- CP-element group 70: 	123 
    -- CP-element group 70: 	124 
    -- CP-element group 70:  members (30) 
      -- CP-element group 70: 	 branch_block_stmt_316/merge_stmt_753__exit__
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794__entry__
      -- CP-element group 70: 	 branch_block_stmt_316/if_stmt_532_if_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_316/if_stmt_532_if_link/if_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_316/forx_xcond119x_xpreheader_bbx_xnph294
      -- CP-element group 70: 	 branch_block_stmt_316/forx_xcond119x_xpreheader_bbx_xnph294_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_update_start_
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_update_start_
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_update_start_
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_316/merge_stmt_753_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_316/merge_stmt_753_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_316/merge_stmt_753_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_316/merge_stmt_753_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_316/forx_xcond119x_xpreheader_bbx_xnph294_PhiReq/$exit
      -- 
    if_choice_transition_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_532_branch_ack_1, ack => zeropad_CP_920_elements(70)); -- 
    rr_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(70), ack => type_cast_756_inst_req_0); -- 
    cr_1854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(70), ack => type_cast_756_inst_req_1); -- 
    rr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(70), ack => type_cast_760_inst_req_0); -- 
    cr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(70), ack => type_cast_760_inst_req_1); -- 
    rr_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(70), ack => type_cast_769_inst_req_0); -- 
    cr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(70), ack => type_cast_769_inst_req_1); -- 
    -- CP-element group 71:  transition  place  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	243 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	256 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_316/if_stmt_532_else_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_316/if_stmt_532_else_link/else_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_316/forx_xcond119x_xpreheader_forx_xend131
      -- CP-element group 71: 	 branch_block_stmt_316/forx_xcond119x_xpreheader_forx_xend131_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_316/forx_xcond119x_xpreheader_forx_xend131_PhiReq/$entry
      -- 
    else_choice_transition_1449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_532_branch_ack_0, ack => zeropad_CP_920_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	68 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_Sample/ra
      -- 
    ra_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_0, ack => zeropad_CP_920_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	68 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	78 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_541_Update/ca
      -- 
    ca_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_1, ack => zeropad_CP_920_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	68 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_Sample/ra
      -- 
    ra_1477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_545_inst_ack_0, ack => zeropad_CP_920_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	68 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_545_Update/ca
      -- 
    ca_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_545_inst_ack_1, ack => zeropad_CP_920_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	68 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_Sample/ra
      -- 
    ra_1491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_554_inst_ack_0, ack => zeropad_CP_920_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	68 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/type_cast_554_Update/ca
      -- 
    ca_1496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_554_inst_ack_1, ack => zeropad_CP_920_elements(77)); -- 
    -- CP-element group 78:  join  transition  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	73 
    -- CP-element group 78: 	75 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	244 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579__exit__
      -- CP-element group 78: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody
      -- CP-element group 78: 	 branch_block_stmt_316/assign_stmt_542_to_assign_stmt_579/$exit
      -- CP-element group 78: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/$entry
      -- CP-element group 78: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody_PhiReq/phi_stmt_582/$entry
      -- CP-element group 78: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody_PhiReq/$entry
      -- 
    zeropad_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(73) & zeropad_CP_920_elements(75) & zeropad_CP_920_elements(77);
      gj_zeropad_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	249 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	118 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_sample_complete
      -- CP-element group 79: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_Sample/ack
      -- 
    ack_1525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_596_index_offset_ack_0, ack => zeropad_CP_920_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	249 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (11) 
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_root_address_calculated
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_offset_calculated
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_Update/ack
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_base_plus_offset/$entry
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_base_plus_offset/$exit
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_base_plus_offset/sum_rename_req
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_base_plus_offset/sum_rename_ack
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_request/$entry
      -- CP-element group 80: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_request/req
      -- 
    ack_1530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_596_index_offset_ack_1, ack => zeropad_CP_920_elements(80)); -- 
    req_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(80), ack => addr_of_597_final_reg_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_request/$exit
      -- CP-element group 81: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_request/ack
      -- 
    ack_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_597_final_reg_ack_0, ack => zeropad_CP_920_elements(81)); -- 
    -- CP-element group 82:  fork  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	249 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	115 
    -- CP-element group 82:  members (19) 
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_complete/$exit
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_complete/ack
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_address_calculated
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_word_address_calculated
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_root_address_calculated
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_address_resized
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_addr_resize/$entry
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_addr_resize/$exit
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_addr_resize/base_resize_req
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_addr_resize/base_resize_ack
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_plus_offset/$entry
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_plus_offset/$exit
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_plus_offset/sum_rename_req
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_base_plus_offset/sum_rename_ack
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_word_addrgen/$entry
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_word_addrgen/$exit
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_word_addrgen/root_register_req
      -- CP-element group 82: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_word_addrgen/root_register_ack
      -- 
    ack_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_597_final_reg_ack_1, ack => zeropad_CP_920_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	249 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_update_start_
      -- CP-element group 83: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_Update/cr
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_600_inst_ack_0, ack => zeropad_CP_920_elements(83)); -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(83), ack => RPIPE_Zeropad_input_pipe_600_inst_req_1); -- 
    -- CP-element group 84:  fork  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	87 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_Sample/rr
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_600_inst_ack_1, ack => zeropad_CP_920_elements(84)); -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(84), ack => RPIPE_Zeropad_input_pipe_613_inst_req_0); -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(84), ack => type_cast_604_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_Sample/ra
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_604_inst_ack_0, ack => zeropad_CP_920_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	249 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	115 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_Update/ca
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_604_inst_ack_1, ack => zeropad_CP_920_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	84 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_update_start_
      -- CP-element group 87: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_Update/cr
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_613_inst_ack_0, ack => zeropad_CP_920_elements(87)); -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(87), ack => RPIPE_Zeropad_input_pipe_613_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	91 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_613_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_Sample/rr
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_613_inst_ack_1, ack => zeropad_CP_920_elements(88)); -- 
    rr_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(88), ack => type_cast_617_inst_req_0); -- 
    rr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(88), ack => RPIPE_Zeropad_input_pipe_631_inst_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_Sample/ra
      -- 
    ra_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_617_inst_ack_0, ack => zeropad_CP_920_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	249 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	115 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_Update/ca
      -- 
    ca_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_617_inst_ack_1, ack => zeropad_CP_920_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	88 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_update_start_
      -- CP-element group 91: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_Update/cr
      -- 
    ra_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_631_inst_ack_0, ack => zeropad_CP_920_elements(91)); -- 
    cr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(91), ack => RPIPE_Zeropad_input_pipe_631_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	95 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_631_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_Sample/rr
      -- 
    ca_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_631_inst_ack_1, ack => zeropad_CP_920_elements(92)); -- 
    rr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(92), ack => RPIPE_Zeropad_input_pipe_649_inst_req_0); -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(92), ack => type_cast_635_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_Sample/ra
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_635_inst_ack_0, ack => zeropad_CP_920_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	249 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	115 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_Update/ca
      -- 
    ca_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_635_inst_ack_1, ack => zeropad_CP_920_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_update_start_
      -- CP-element group 95: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_Update/cr
      -- 
    ra_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_649_inst_ack_0, ack => zeropad_CP_920_elements(95)); -- 
    cr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(95), ack => RPIPE_Zeropad_input_pipe_649_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	99 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_649_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_Sample/rr
      -- 
    ca_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_649_inst_ack_1, ack => zeropad_CP_920_elements(96)); -- 
    rr_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(96), ack => type_cast_653_inst_req_0); -- 
    rr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(96), ack => RPIPE_Zeropad_input_pipe_667_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_Sample/ra
      -- 
    ra_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_653_inst_ack_0, ack => zeropad_CP_920_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	249 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	115 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_Update/ca
      -- 
    ca_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_653_inst_ack_1, ack => zeropad_CP_920_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_update_start_
      -- CP-element group 99: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_Update/cr
      -- 
    ra_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_667_inst_ack_0, ack => zeropad_CP_920_elements(99)); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(99), ack => RPIPE_Zeropad_input_pipe_667_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_667_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_Sample/rr
      -- 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_667_inst_ack_1, ack => zeropad_CP_920_elements(100)); -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(100), ack => type_cast_671_inst_req_0); -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(100), ack => RPIPE_Zeropad_input_pipe_685_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_Sample/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_671_inst_ack_0, ack => zeropad_CP_920_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	249 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	115 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_Update/ca
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_671_inst_ack_1, ack => zeropad_CP_920_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_update_start_
      -- CP-element group 103: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_Update/cr
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_685_inst_ack_0, ack => zeropad_CP_920_elements(103)); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(103), ack => RPIPE_Zeropad_input_pipe_685_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_685_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_Sample/rr
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_685_inst_ack_1, ack => zeropad_CP_920_elements(104)); -- 
    rr_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(104), ack => type_cast_689_inst_req_0); -- 
    rr_1721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(104), ack => RPIPE_Zeropad_input_pipe_703_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_Sample/ra
      -- 
    ra_1708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_689_inst_ack_0, ack => zeropad_CP_920_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	249 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	115 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_Update/ca
      -- 
    ca_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_689_inst_ack_1, ack => zeropad_CP_920_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_update_start_
      -- CP-element group 107: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_Update/cr
      -- 
    ra_1722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_703_inst_ack_0, ack => zeropad_CP_920_elements(107)); -- 
    cr_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(107), ack => RPIPE_Zeropad_input_pipe_703_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	111 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_703_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_Sample/rr
      -- 
    ca_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_703_inst_ack_1, ack => zeropad_CP_920_elements(108)); -- 
    rr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(108), ack => RPIPE_Zeropad_input_pipe_721_inst_req_0); -- 
    rr_1735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(108), ack => type_cast_707_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_Sample/ra
      -- 
    ra_1736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_707_inst_ack_0, ack => zeropad_CP_920_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	249 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	115 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_Update/ca
      -- 
    ca_1741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_707_inst_ack_1, ack => zeropad_CP_920_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_update_start_
      -- CP-element group 111: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_Update/cr
      -- 
    ra_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_721_inst_ack_0, ack => zeropad_CP_920_elements(111)); -- 
    cr_1754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(111), ack => RPIPE_Zeropad_input_pipe_721_inst_req_1); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_721_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_Sample/rr
      -- 
    ca_1755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_721_inst_ack_1, ack => zeropad_CP_920_elements(112)); -- 
    rr_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(112), ack => type_cast_725_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_Sample/ra
      -- 
    ra_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_725_inst_ack_0, ack => zeropad_CP_920_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	249 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_Update/ca
      -- 
    ca_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_725_inst_ack_1, ack => zeropad_CP_920_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	86 
    -- CP-element group 115: 	94 
    -- CP-element group 115: 	82 
    -- CP-element group 115: 	90 
    -- CP-element group 115: 	114 
    -- CP-element group 115: 	106 
    -- CP-element group 115: 	110 
    -- CP-element group 115: 	98 
    -- CP-element group 115: 	102 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (9) 
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/ptr_deref_733_Split/$entry
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/ptr_deref_733_Split/$exit
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/ptr_deref_733_Split/split_req
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/ptr_deref_733_Split/split_ack
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/word_access_start/$entry
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/word_access_start/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/word_access_start/word_0/rr
      -- 
    rr_1807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(115), ack => ptr_deref_733_store_0_req_0); -- 
    zeropad_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(86) & zeropad_CP_920_elements(94) & zeropad_CP_920_elements(82) & zeropad_CP_920_elements(90) & zeropad_CP_920_elements(114) & zeropad_CP_920_elements(106) & zeropad_CP_920_elements(110) & zeropad_CP_920_elements(98) & zeropad_CP_920_elements(102);
      gj_zeropad_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/word_access_start/$exit
      -- CP-element group 116: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/word_access_start/word_0/$exit
      -- CP-element group 116: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Sample/word_access_start/word_0/ra
      -- 
    ra_1808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_733_store_0_ack_0, ack => zeropad_CP_920_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	249 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Update/word_access_complete/$exit
      -- CP-element group 117: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Update/word_access_complete/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Update/word_access_complete/word_0/ca
      -- 
    ca_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_733_store_0_ack_1, ack => zeropad_CP_920_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	79 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746__exit__
      -- CP-element group 118: 	 branch_block_stmt_316/if_stmt_747__entry__
      -- CP-element group 118: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/$exit
      -- CP-element group 118: 	 branch_block_stmt_316/if_stmt_747_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_316/if_stmt_747_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_316/if_stmt_747_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_316/if_stmt_747_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_316/R_exitcond24_748_place
      -- CP-element group 118: 	 branch_block_stmt_316/if_stmt_747_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_316/if_stmt_747_else_link/$entry
      -- 
    branch_req_1827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(118), ack => if_stmt_747_branch_req_0); -- 
    zeropad_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(79) & zeropad_CP_920_elements(117);
      gj_zeropad_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  transition  place  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	243 
    -- CP-element group 119:  members (13) 
      -- CP-element group 119: 	 branch_block_stmt_316/merge_stmt_523__exit__
      -- CP-element group 119: 	 branch_block_stmt_316/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader
      -- CP-element group 119: 	 branch_block_stmt_316/if_stmt_747_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_316/if_stmt_747_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_316/forx_xbody_forx_xcond119x_xpreheaderx_xloopexit
      -- CP-element group 119: 	 branch_block_stmt_316/forx_xbody_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_316/forx_xbody_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_316/merge_stmt_523_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_316/merge_stmt_523_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_316/merge_stmt_523_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_316/merge_stmt_523_PhiAck/dummy
      -- CP-element group 119: 	 branch_block_stmt_316/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_316/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_747_branch_ack_1, ack => zeropad_CP_920_elements(119)); -- 
    -- CP-element group 120:  fork  transition  place  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	245 
    -- CP-element group 120: 	246 
    -- CP-element group 120:  members (12) 
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/$entry
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/$entry
      -- CP-element group 120: 	 branch_block_stmt_316/if_stmt_747_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_316/if_stmt_747_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/Update/cr
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/$entry
      -- CP-element group 120: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/$entry
      -- 
    else_choice_transition_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_747_branch_ack_0, ack => zeropad_CP_920_elements(120)); -- 
    cr_2780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(120), ack => type_cast_588_inst_req_1); -- 
    rr_2775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(120), ack => type_cast_588_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	70 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_Sample/ra
      -- 
    ra_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_756_inst_ack_0, ack => zeropad_CP_920_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	70 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	127 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_756_Update/ca
      -- 
    ca_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_756_inst_ack_1, ack => zeropad_CP_920_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	70 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_Sample/ra
      -- 
    ra_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_760_inst_ack_0, ack => zeropad_CP_920_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	70 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_760_Update/ca
      -- 
    ca_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_760_inst_ack_1, ack => zeropad_CP_920_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	70 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_Sample/ra
      -- 
    ra_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_0, ack => zeropad_CP_920_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	70 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/type_cast_769_Update/ca
      -- 
    ca_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_1, ack => zeropad_CP_920_elements(126)); -- 
    -- CP-element group 127:  join  transition  place  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: 	122 
    -- CP-element group 127: 	124 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	250 
    -- CP-element group 127:  members (6) 
      -- CP-element group 127: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794__exit__
      -- CP-element group 127: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125
      -- CP-element group 127: 	 branch_block_stmt_316/assign_stmt_757_to_assign_stmt_794/$exit
      -- CP-element group 127: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125_PhiReq/phi_stmt_797/$entry
      -- CP-element group 127: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125_PhiReq/$entry
      -- 
    zeropad_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(126) & zeropad_CP_920_elements(122) & zeropad_CP_920_elements(124);
      gj_zeropad_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	255 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	134 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_sample_complete
      -- CP-element group 128: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_Sample/ack
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_811_index_offset_ack_0, ack => zeropad_CP_920_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	255 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (11) 
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_request/req
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_request/$entry
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_base_plus_offset/sum_rename_ack
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_root_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_offset_calculated
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_Update/ack
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_base_plus_offset/$entry
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_base_plus_offset/$exit
      -- CP-element group 129: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_base_plus_offset/sum_rename_req
      -- 
    ack_1917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_811_index_offset_ack_1, ack => zeropad_CP_920_elements(129)); -- 
    req_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(129), ack => addr_of_812_final_reg_req_0); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_request/ack
      -- CP-element group 130: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_request/$exit
      -- CP-element group 130: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_sample_completed_
      -- 
    ack_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_812_final_reg_ack_0, ack => zeropad_CP_920_elements(130)); -- 
    -- CP-element group 131:  join  fork  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	255 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (28) 
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_complete/ack
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_complete/$exit
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_word_addrgen/root_register_ack
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_address_calculated
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_word_address_calculated
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_root_address_calculated
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_address_resized
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_addr_resize/$entry
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_addr_resize/$exit
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_addr_resize/base_resize_req
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_addr_resize/base_resize_ack
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_plus_offset/$entry
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_plus_offset/$exit
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_plus_offset/sum_rename_req
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_base_plus_offset/sum_rename_ack
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/ptr_deref_815_Split/$entry
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/ptr_deref_815_Split/$exit
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_word_addrgen/$entry
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_word_addrgen/$exit
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/word_access_start/word_0/rr
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/word_access_start/word_0/$entry
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/word_access_start/$entry
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_word_addrgen/root_register_req
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/ptr_deref_815_Split/split_ack
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/ptr_deref_815_Split/split_req
      -- CP-element group 131: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_update_completed_
      -- 
    ack_1932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_812_final_reg_ack_1, ack => zeropad_CP_920_elements(131)); -- 
    rr_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(131), ack => ptr_deref_815_store_0_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/word_access_start/word_0/ra
      -- CP-element group 132: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/word_access_start/word_0/$exit
      -- CP-element group 132: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Sample/word_access_start/$exit
      -- 
    ra_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_815_store_0_ack_0, ack => zeropad_CP_920_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	255 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Update/word_access_complete/word_0/ca
      -- CP-element group 133: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Update/word_access_complete/word_0/$exit
      -- CP-element group 133: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Update/word_access_complete/$exit
      -- CP-element group 133: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Update/$exit
      -- 
    ca_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_815_store_0_ack_1, ack => zeropad_CP_920_elements(133)); -- 
    -- CP-element group 134:  branch  join  transition  place  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	128 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (10) 
      -- CP-element group 134: 	 branch_block_stmt_316/if_stmt_830_dead_link/$entry
      -- CP-element group 134: 	 branch_block_stmt_316/if_stmt_830_eval_test/branch_req
      -- CP-element group 134: 	 branch_block_stmt_316/if_stmt_830_else_link/$entry
      -- CP-element group 134: 	 branch_block_stmt_316/if_stmt_830_eval_test/$entry
      -- CP-element group 134: 	 branch_block_stmt_316/if_stmt_830_eval_test/$exit
      -- CP-element group 134: 	 branch_block_stmt_316/if_stmt_830_if_link/$entry
      -- CP-element group 134: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829__exit__
      -- CP-element group 134: 	 branch_block_stmt_316/if_stmt_830__entry__
      -- CP-element group 134: 	 branch_block_stmt_316/R_exitcond_831_place
      -- CP-element group 134: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/$exit
      -- 
    branch_req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(134), ack => if_stmt_830_branch_req_0); -- 
    zeropad_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(128) & zeropad_CP_920_elements(133);
      gj_zeropad_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  merge  transition  place  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	256 
    -- CP-element group 135:  members (13) 
      -- CP-element group 135: 	 branch_block_stmt_316/if_stmt_830_if_link/$exit
      -- CP-element group 135: 	 branch_block_stmt_316/if_stmt_830_if_link/if_choice_transition
      -- CP-element group 135: 	 branch_block_stmt_316/merge_stmt_836__exit__
      -- CP-element group 135: 	 branch_block_stmt_316/forx_xend131x_xloopexit_forx_xend131
      -- CP-element group 135: 	 branch_block_stmt_316/forx_xbody125_forx_xend131x_xloopexit
      -- CP-element group 135: 	 branch_block_stmt_316/forx_xbody125_forx_xend131x_xloopexit_PhiReq/$entry
      -- CP-element group 135: 	 branch_block_stmt_316/forx_xbody125_forx_xend131x_xloopexit_PhiReq/$exit
      -- CP-element group 135: 	 branch_block_stmt_316/merge_stmt_836_PhiReqMerge
      -- CP-element group 135: 	 branch_block_stmt_316/forx_xend131x_xloopexit_forx_xend131_PhiReq/$exit
      -- CP-element group 135: 	 branch_block_stmt_316/forx_xend131x_xloopexit_forx_xend131_PhiReq/$entry
      -- CP-element group 135: 	 branch_block_stmt_316/merge_stmt_836_PhiAck/dummy
      -- CP-element group 135: 	 branch_block_stmt_316/merge_stmt_836_PhiAck/$exit
      -- CP-element group 135: 	 branch_block_stmt_316/merge_stmt_836_PhiAck/$entry
      -- 
    if_choice_transition_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_830_branch_ack_1, ack => zeropad_CP_920_elements(135)); -- 
    -- CP-element group 136:  fork  transition  place  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	251 
    -- CP-element group 136: 	252 
    -- CP-element group 136:  members (12) 
      -- CP-element group 136: 	 branch_block_stmt_316/if_stmt_830_else_link/$exit
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/$entry
      -- CP-element group 136: 	 branch_block_stmt_316/if_stmt_830_else_link/else_choice_transition
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/$entry
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/$entry
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/$entry
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/$entry
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/Sample/rr
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_830_branch_ack_0, ack => zeropad_CP_920_elements(136)); -- 
    rr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(136), ack => type_cast_803_inst_req_0); -- 
    cr_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(136), ack => type_cast_803_inst_req_1); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	256 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_Sample/cra
      -- 
    cra_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_841_call_ack_0, ack => zeropad_CP_920_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	256 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_Update/cca
      -- CP-element group 138: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_Sample/rr
      -- 
    cca_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_841_call_ack_1, ack => zeropad_CP_920_elements(138)); -- 
    rr_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(138), ack => type_cast_846_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_Sample/ra
      -- 
    ra_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_846_inst_ack_0, ack => zeropad_CP_920_elements(139)); -- 
    -- CP-element group 140:  fork  transition  place  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	256 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (13) 
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/$exit
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847__exit__
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_859__entry__
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_Update/ccr
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_Sample/crr
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_update_start_
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_859/$entry
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_Update/$exit
      -- 
    ca_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_846_inst_ack_1, ack => zeropad_CP_920_elements(140)); -- 
    ccr_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(140), ack => call_stmt_859_call_req_1); -- 
    crr_2043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(140), ack => call_stmt_859_call_req_0); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_Sample/cra
      -- CP-element group 141: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_sample_completed_
      -- 
    cra_2044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_859_call_ack_0, ack => zeropad_CP_920_elements(141)); -- 
    -- CP-element group 142:  fork  transition  place  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	144 
    -- CP-element group 142: 	146 
    -- CP-element group 142: 	148 
    -- CP-element group 142: 	150 
    -- CP-element group 142: 	152 
    -- CP-element group 142: 	154 
    -- CP-element group 142: 	156 
    -- CP-element group 142: 	158 
    -- CP-element group 142: 	160 
    -- CP-element group 142: 	162 
    -- CP-element group 142:  members (40) 
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_Update/ccr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_Sample/crr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_859__exit__
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970__entry__
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_Update/cca
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_859/call_stmt_859_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_859/$exit
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_update_start_
      -- CP-element group 142: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_Update/cr
      -- 
    cca_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_859_call_ack_1, ack => zeropad_CP_920_elements(142)); -- 
    cr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_945_inst_req_1); -- 
    cr_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_915_inst_req_1); -- 
    ccr_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => call_stmt_862_call_req_1); -- 
    crr_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => call_stmt_862_call_req_0); -- 
    cr_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_925_inst_req_1); -- 
    cr_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_866_inst_req_1); -- 
    cr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_875_inst_req_1); -- 
    cr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_885_inst_req_1); -- 
    cr_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_905_inst_req_1); -- 
    cr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_935_inst_req_1); -- 
    cr_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(142), ack => type_cast_895_inst_req_1); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_Sample/cra
      -- CP-element group 143: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_sample_completed_
      -- 
    cra_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_862_call_ack_0, ack => zeropad_CP_920_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (6) 
      -- CP-element group 144: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_Update/cca
      -- CP-element group 144: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/call_stmt_862_update_completed_
      -- 
    cca_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_862_call_ack_1, ack => zeropad_CP_920_elements(144)); -- 
    rr_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(144), ack => type_cast_866_inst_req_0); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_Sample/ra
      -- 
    ra_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_866_inst_ack_0, ack => zeropad_CP_920_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	142 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146: 	151 
    -- CP-element group 146: 	153 
    -- CP-element group 146: 	155 
    -- CP-element group 146: 	157 
    -- CP-element group 146: 	159 
    -- CP-element group 146: 	161 
    -- CP-element group 146:  members (27) 
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_866_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_sample_start_
      -- 
    ca_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_866_inst_ack_1, ack => zeropad_CP_920_elements(146)); -- 
    rr_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(146), ack => type_cast_875_inst_req_0); -- 
    rr_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(146), ack => type_cast_885_inst_req_0); -- 
    rr_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(146), ack => type_cast_895_inst_req_0); -- 
    rr_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(146), ack => type_cast_905_inst_req_0); -- 
    rr_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(146), ack => type_cast_915_inst_req_0); -- 
    rr_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(146), ack => type_cast_925_inst_req_0); -- 
    rr_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(146), ack => type_cast_935_inst_req_0); -- 
    rr_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(146), ack => type_cast_945_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_Sample/ra
      -- 
    ra_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_875_inst_ack_0, ack => zeropad_CP_920_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	142 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	183 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_875_Update/ca
      -- 
    ca_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_875_inst_ack_1, ack => zeropad_CP_920_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_Sample/ra
      -- 
    ra_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_885_inst_ack_0, ack => zeropad_CP_920_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	142 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	180 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_885_Update/$exit
      -- 
    ca_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_885_inst_ack_1, ack => zeropad_CP_920_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	146 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_sample_completed_
      -- 
    ra_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_895_inst_ack_0, ack => zeropad_CP_920_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	142 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	177 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_895_Update/ca
      -- 
    ca_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_895_inst_ack_1, ack => zeropad_CP_920_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	146 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_sample_completed_
      -- 
    ra_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_0, ack => zeropad_CP_920_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	142 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	174 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_905_update_completed_
      -- 
    ca_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_1, ack => zeropad_CP_920_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	146 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_sample_completed_
      -- 
    ra_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_0, ack => zeropad_CP_920_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	142 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	171 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_915_update_completed_
      -- 
    ca_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_1, ack => zeropad_CP_920_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	146 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_Sample/ra
      -- 
    ra_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_925_inst_ack_0, ack => zeropad_CP_920_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	142 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	168 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_925_Update/ca
      -- 
    ca_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_925_inst_ack_1, ack => zeropad_CP_920_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	146 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_Sample/ra
      -- 
    ra_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_935_inst_ack_0, ack => zeropad_CP_920_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	142 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	165 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_935_Update/ca
      -- 
    ca_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_935_inst_ack_1, ack => zeropad_CP_920_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	146 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_Sample/ra
      -- CP-element group 161: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_sample_completed_
      -- 
    ra_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_945_inst_ack_0, ack => zeropad_CP_920_elements(161)); -- 
    -- CP-element group 162:  transition  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	142 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (6) 
      -- CP-element group 162: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_Update/ca
      -- CP-element group 162: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/type_cast_945_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_Sample/req
      -- 
    ca_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_945_inst_ack_1, ack => zeropad_CP_920_elements(162)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(162), ack => WPIPE_Zeropad_output_pipe_947_inst_req_0); -- 
    -- CP-element group 163:  transition  input  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (6) 
      -- CP-element group 163: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_Update/req
      -- CP-element group 163: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_update_start_
      -- CP-element group 163: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_Sample/ack
      -- CP-element group 163: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_Sample/$exit
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_947_inst_ack_0, ack => zeropad_CP_920_elements(163)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(163), ack => WPIPE_Zeropad_output_pipe_947_inst_req_1); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_Update/ack
      -- CP-element group 164: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_947_update_completed_
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_947_inst_ack_1, ack => zeropad_CP_920_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	160 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_Sample/req
      -- CP-element group 165: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_Sample/$entry
      -- 
    req_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(165), ack => WPIPE_Zeropad_output_pipe_950_inst_req_0); -- 
    zeropad_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(160) & zeropad_CP_920_elements(164);
      gj_zeropad_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (6) 
      -- CP-element group 166: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_update_start_
      -- CP-element group 166: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_Update/req
      -- CP-element group 166: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_Sample/ack
      -- CP-element group 166: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_Sample/$exit
      -- 
    ack_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_950_inst_ack_0, ack => zeropad_CP_920_elements(166)); -- 
    req_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(166), ack => WPIPE_Zeropad_output_pipe_950_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_Update/ack
      -- CP-element group 167: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_950_update_completed_
      -- 
    ack_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_950_inst_ack_1, ack => zeropad_CP_920_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	158 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_Sample/req
      -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(168), ack => WPIPE_Zeropad_output_pipe_953_inst_req_0); -- 
    zeropad_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(158) & zeropad_CP_920_elements(167);
      gj_zeropad_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (6) 
      -- CP-element group 169: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_update_start_
      -- CP-element group 169: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_Update/req
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_953_inst_ack_0, ack => zeropad_CP_920_elements(169)); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(169), ack => WPIPE_Zeropad_output_pipe_953_inst_req_1); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_953_Update/ack
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_953_inst_ack_1, ack => zeropad_CP_920_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	156 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_Sample/req
      -- CP-element group 171: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_sample_start_
      -- 
    req_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(171), ack => WPIPE_Zeropad_output_pipe_956_inst_req_0); -- 
    zeropad_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(156) & zeropad_CP_920_elements(170);
      gj_zeropad_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_Update/req
      -- CP-element group 172: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_Sample/ack
      -- CP-element group 172: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_update_start_
      -- CP-element group 172: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_sample_completed_
      -- 
    ack_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_956_inst_ack_0, ack => zeropad_CP_920_elements(172)); -- 
    req_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(172), ack => WPIPE_Zeropad_output_pipe_956_inst_req_1); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_Update/ack
      -- CP-element group 173: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_956_update_completed_
      -- 
    ack_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_956_inst_ack_1, ack => zeropad_CP_920_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	154 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_Sample/req
      -- CP-element group 174: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_sample_start_
      -- 
    req_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(174), ack => WPIPE_Zeropad_output_pipe_959_inst_req_0); -- 
    zeropad_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(154) & zeropad_CP_920_elements(173);
      gj_zeropad_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_Sample/ack
      -- CP-element group 175: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_update_start_
      -- CP-element group 175: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_Update/req
      -- CP-element group 175: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_Update/$entry
      -- 
    ack_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_959_inst_ack_0, ack => zeropad_CP_920_elements(175)); -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(175), ack => WPIPE_Zeropad_output_pipe_959_inst_req_1); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_Update/ack
      -- CP-element group 176: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_959_Update/$exit
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_959_inst_ack_1, ack => zeropad_CP_920_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	152 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_Sample/req
      -- CP-element group 177: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_sample_start_
      -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(177), ack => WPIPE_Zeropad_output_pipe_962_inst_req_0); -- 
    zeropad_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(152) & zeropad_CP_920_elements(176);
      gj_zeropad_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (6) 
      -- CP-element group 178: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_Sample/ack
      -- CP-element group 178: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_Update/req
      -- CP-element group 178: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_update_start_
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_962_inst_ack_0, ack => zeropad_CP_920_elements(178)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(178), ack => WPIPE_Zeropad_output_pipe_962_inst_req_1); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_Update/ack
      -- CP-element group 179: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_962_update_completed_
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_962_inst_ack_1, ack => zeropad_CP_920_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	150 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_Sample/req
      -- CP-element group 180: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_Sample/$entry
      -- 
    req_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(180), ack => WPIPE_Zeropad_output_pipe_965_inst_req_0); -- 
    zeropad_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(150) & zeropad_CP_920_elements(179);
      gj_zeropad_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_Sample/ack
      -- CP-element group 181: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_Update/req
      -- CP-element group 181: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_update_start_
      -- 
    ack_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_965_inst_ack_0, ack => zeropad_CP_920_elements(181)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(181), ack => WPIPE_Zeropad_output_pipe_965_inst_req_1); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_965_Update/ack
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_965_inst_ack_1, ack => zeropad_CP_920_elements(182)); -- 
    -- CP-element group 183:  join  transition  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	148 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_Sample/req
      -- 
    req_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(183), ack => WPIPE_Zeropad_output_pipe_968_inst_req_0); -- 
    zeropad_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(148) & zeropad_CP_920_elements(182);
      gj_zeropad_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (6) 
      -- CP-element group 184: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_update_start_
      -- CP-element group 184: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_Sample/ack
      -- CP-element group 184: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_Update/req
      -- 
    ack_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_968_inst_ack_0, ack => zeropad_CP_920_elements(184)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(184), ack => WPIPE_Zeropad_output_pipe_968_inst_req_1); -- 
    -- CP-element group 185:  branch  transition  place  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (13) 
      -- CP-element group 185: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970__exit__
      -- CP-element group 185: 	 branch_block_stmt_316/if_stmt_972__entry__
      -- CP-element group 185: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/$exit
      -- CP-element group 185: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_316/call_stmt_862_to_assign_stmt_970/WPIPE_Zeropad_output_pipe_968_Update/ack
      -- CP-element group 185: 	 branch_block_stmt_316/if_stmt_972_dead_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_316/if_stmt_972_eval_test/$entry
      -- CP-element group 185: 	 branch_block_stmt_316/if_stmt_972_eval_test/$exit
      -- CP-element group 185: 	 branch_block_stmt_316/if_stmt_972_eval_test/branch_req
      -- CP-element group 185: 	 branch_block_stmt_316/R_cmp123292_973_place
      -- CP-element group 185: 	 branch_block_stmt_316/if_stmt_972_if_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_316/if_stmt_972_else_link/$entry
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_968_inst_ack_1, ack => zeropad_CP_920_elements(185)); -- 
    branch_req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(185), ack => if_stmt_972_branch_req_0); -- 
    -- CP-element group 186:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: 	189 
    -- CP-element group 186: 	190 
    -- CP-element group 186: 	191 
    -- CP-element group 186: 	192 
    -- CP-element group 186: 	193 
    -- CP-element group 186:  members (30) 
      -- CP-element group 186: 	 branch_block_stmt_316/merge_stmt_978_PhiReqMerge
      -- CP-element group 186: 	 branch_block_stmt_316/merge_stmt_978__exit__
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019__entry__
      -- CP-element group 186: 	 branch_block_stmt_316/if_stmt_972_if_link/$exit
      -- CP-element group 186: 	 branch_block_stmt_316/if_stmt_972_if_link/if_choice_transition
      -- CP-element group 186: 	 branch_block_stmt_316/forx_xend131_bbx_xnph
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/$entry
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_update_start_
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_update_start_
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_update_start_
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_316/merge_stmt_978_PhiAck/dummy
      -- CP-element group 186: 	 branch_block_stmt_316/merge_stmt_978_PhiAck/$exit
      -- CP-element group 186: 	 branch_block_stmt_316/merge_stmt_978_PhiAck/$entry
      -- CP-element group 186: 	 branch_block_stmt_316/forx_xend131_bbx_xnph_PhiReq/$exit
      -- CP-element group 186: 	 branch_block_stmt_316/forx_xend131_bbx_xnph_PhiReq/$entry
      -- 
    if_choice_transition_2317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_972_branch_ack_1, ack => zeropad_CP_920_elements(186)); -- 
    rr_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(186), ack => type_cast_981_inst_req_0); -- 
    cr_2339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(186), ack => type_cast_981_inst_req_1); -- 
    rr_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(186), ack => type_cast_985_inst_req_0); -- 
    cr_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(186), ack => type_cast_985_inst_req_1); -- 
    rr_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(186), ack => type_cast_994_inst_req_0); -- 
    cr_2367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(186), ack => type_cast_994_inst_req_1); -- 
    -- CP-element group 187:  transition  place  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	263 
    -- CP-element group 187:  members (5) 
      -- CP-element group 187: 	 branch_block_stmt_316/forx_xend131_forx_xend287_PhiReq/$entry
      -- CP-element group 187: 	 branch_block_stmt_316/forx_xend131_forx_xend287_PhiReq/$exit
      -- CP-element group 187: 	 branch_block_stmt_316/if_stmt_972_else_link/$exit
      -- CP-element group 187: 	 branch_block_stmt_316/if_stmt_972_else_link/else_choice_transition
      -- CP-element group 187: 	 branch_block_stmt_316/forx_xend131_forx_xend287
      -- 
    else_choice_transition_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_972_branch_ack_0, ack => zeropad_CP_920_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_Sample/ra
      -- 
    ra_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_981_inst_ack_0, ack => zeropad_CP_920_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	194 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_981_Update/ca
      -- 
    ca_2340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_981_inst_ack_1, ack => zeropad_CP_920_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	186 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_Sample/ra
      -- 
    ra_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_985_inst_ack_0, ack => zeropad_CP_920_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	186 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	194 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_985_Update/ca
      -- 
    ca_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_985_inst_ack_1, ack => zeropad_CP_920_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	186 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_Sample/ra
      -- 
    ra_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_994_inst_ack_0, ack => zeropad_CP_920_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	186 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/type_cast_994_Update/ca
      -- 
    ca_2368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_994_inst_ack_1, ack => zeropad_CP_920_elements(193)); -- 
    -- CP-element group 194:  join  transition  place  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	189 
    -- CP-element group 194: 	191 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	257 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019__exit__
      -- CP-element group 194: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215
      -- CP-element group 194: 	 branch_block_stmt_316/assign_stmt_982_to_assign_stmt_1019/$exit
      -- CP-element group 194: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/$entry
      -- CP-element group 194: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215_PhiReq/phi_stmt_1022/$entry
      -- CP-element group 194: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215_PhiReq/$entry
      -- 
    zeropad_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(189) & zeropad_CP_920_elements(191) & zeropad_CP_920_elements(193);
      gj_zeropad_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	262 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	240 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_sample_complete
      -- CP-element group 195: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_Sample/ack
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1036_index_offset_ack_0, ack => zeropad_CP_920_elements(195)); -- 
    -- CP-element group 196:  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	262 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (11) 
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_root_address_calculated
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_offset_calculated
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_Update/ack
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_base_plus_offset/$entry
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_base_plus_offset/$exit
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_base_plus_offset/sum_rename_req
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_base_plus_offset/sum_rename_ack
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_request/$entry
      -- CP-element group 196: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_request/req
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1036_index_offset_ack_1, ack => zeropad_CP_920_elements(196)); -- 
    req_2411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(196), ack => addr_of_1037_final_reg_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_request/$exit
      -- CP-element group 197: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_request/ack
      -- 
    ack_2412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1037_final_reg_ack_0, ack => zeropad_CP_920_elements(197)); -- 
    -- CP-element group 198:  join  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	262 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (24) 
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_complete/$exit
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_complete/ack
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_address_calculated
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_word_address_calculated
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_root_address_calculated
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_address_resized
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_addr_resize/$entry
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_addr_resize/$exit
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_addr_resize/base_resize_req
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_addr_resize/base_resize_ack
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_plus_offset/$entry
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_plus_offset/$exit
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_plus_offset/sum_rename_req
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_base_plus_offset/sum_rename_ack
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_word_addrgen/$entry
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_word_addrgen/$exit
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_word_addrgen/root_register_req
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_word_addrgen/root_register_ack
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Sample/word_access_start/$entry
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Sample/word_access_start/word_0/$entry
      -- CP-element group 198: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Sample/word_access_start/word_0/rr
      -- 
    ack_2417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1037_final_reg_ack_1, ack => zeropad_CP_920_elements(198)); -- 
    rr_2450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(198), ack => ptr_deref_1041_load_0_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (5) 
      -- CP-element group 199: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Sample/word_access_start/$exit
      -- CP-element group 199: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Sample/word_access_start/word_0/$exit
      -- CP-element group 199: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Sample/word_access_start/word_0/ra
      -- 
    ra_2451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_0_ack_0, ack => zeropad_CP_920_elements(199)); -- 
    -- CP-element group 200:  fork  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	262 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	203 
    -- CP-element group 200: 	205 
    -- CP-element group 200: 	207 
    -- CP-element group 200: 	209 
    -- CP-element group 200: 	211 
    -- CP-element group 200: 	213 
    -- CP-element group 200: 	215 
    -- CP-element group 200:  members (33) 
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/word_access_complete/$exit
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/word_access_complete/word_0/$exit
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/word_access_complete/word_0/ca
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/ptr_deref_1041_Merge/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/ptr_deref_1041_Merge/$exit
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/ptr_deref_1041_Merge/merge_req
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/ptr_deref_1041_Merge/merge_ack
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_Sample/rr
      -- 
    ca_2462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_0_ack_1, ack => zeropad_CP_920_elements(200)); -- 
    rr_2475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(200), ack => type_cast_1045_inst_req_0); -- 
    rr_2489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(200), ack => type_cast_1055_inst_req_0); -- 
    rr_2503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(200), ack => type_cast_1065_inst_req_0); -- 
    rr_2517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(200), ack => type_cast_1075_inst_req_0); -- 
    rr_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(200), ack => type_cast_1085_inst_req_0); -- 
    rr_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(200), ack => type_cast_1095_inst_req_0); -- 
    rr_2559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(200), ack => type_cast_1105_inst_req_0); -- 
    rr_2573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(200), ack => type_cast_1115_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_Sample/ra
      -- 
    ra_2476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1045_inst_ack_0, ack => zeropad_CP_920_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	262 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	237 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_Update/ca
      -- 
    ca_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1045_inst_ack_1, ack => zeropad_CP_920_elements(202)); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	200 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_Sample/ra
      -- 
    ra_2490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_0, ack => zeropad_CP_920_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	262 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	234 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_Update/ca
      -- 
    ca_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_1, ack => zeropad_CP_920_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	200 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_Sample/ra
      -- 
    ra_2504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1065_inst_ack_0, ack => zeropad_CP_920_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	262 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	231 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_Update/ca
      -- 
    ca_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1065_inst_ack_1, ack => zeropad_CP_920_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	200 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_Sample/ra
      -- 
    ra_2518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1075_inst_ack_0, ack => zeropad_CP_920_elements(207)); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	262 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	228 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_Update/ca
      -- 
    ca_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1075_inst_ack_1, ack => zeropad_CP_920_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	200 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_Sample/ra
      -- 
    ra_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_0, ack => zeropad_CP_920_elements(209)); -- 
    -- CP-element group 210:  transition  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	262 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	225 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_Update/ca
      -- 
    ca_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_1, ack => zeropad_CP_920_elements(210)); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	200 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_Sample/ra
      -- 
    ra_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1095_inst_ack_0, ack => zeropad_CP_920_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	262 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	222 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_Update/ca
      -- 
    ca_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1095_inst_ack_1, ack => zeropad_CP_920_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	200 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_Sample/ra
      -- 
    ra_2560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_0, ack => zeropad_CP_920_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	262 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	219 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_Update/ca
      -- 
    ca_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_1, ack => zeropad_CP_920_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	200 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_Sample/ra
      -- 
    ra_2574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1115_inst_ack_0, ack => zeropad_CP_920_elements(215)); -- 
    -- CP-element group 216:  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	262 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_Sample/req
      -- 
    ca_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1115_inst_ack_1, ack => zeropad_CP_920_elements(216)); -- 
    req_2587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(216), ack => WPIPE_Zeropad_output_pipe_1117_inst_req_0); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_update_start_
      -- CP-element group 217: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_Sample/ack
      -- CP-element group 217: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_Update/req
      -- 
    ack_2588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1117_inst_ack_0, ack => zeropad_CP_920_elements(217)); -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(217), ack => WPIPE_Zeropad_output_pipe_1117_inst_req_1); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1117_Update/ack
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1117_inst_ack_1, ack => zeropad_CP_920_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	214 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_Sample/req
      -- 
    req_2601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(219), ack => WPIPE_Zeropad_output_pipe_1120_inst_req_0); -- 
    zeropad_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(214) & zeropad_CP_920_elements(218);
      gj_zeropad_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (6) 
      -- CP-element group 220: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_update_start_
      -- CP-element group 220: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_Sample/ack
      -- CP-element group 220: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_Update/req
      -- 
    ack_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1120_inst_ack_0, ack => zeropad_CP_920_elements(220)); -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(220), ack => WPIPE_Zeropad_output_pipe_1120_inst_req_1); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1120_Update/ack
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1120_inst_ack_1, ack => zeropad_CP_920_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	212 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_Sample/req
      -- 
    req_2615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(222), ack => WPIPE_Zeropad_output_pipe_1123_inst_req_0); -- 
    zeropad_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(212) & zeropad_CP_920_elements(221);
      gj_zeropad_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (6) 
      -- CP-element group 223: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_update_start_
      -- CP-element group 223: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_Update/req
      -- 
    ack_2616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1123_inst_ack_0, ack => zeropad_CP_920_elements(223)); -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(223), ack => WPIPE_Zeropad_output_pipe_1123_inst_req_1); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1123_Update/ack
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1123_inst_ack_1, ack => zeropad_CP_920_elements(224)); -- 
    -- CP-element group 225:  join  transition  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	210 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_Sample/req
      -- 
    req_2629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(225), ack => WPIPE_Zeropad_output_pipe_1126_inst_req_0); -- 
    zeropad_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(210) & zeropad_CP_920_elements(224);
      gj_zeropad_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (6) 
      -- CP-element group 226: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_update_start_
      -- CP-element group 226: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_Sample/ack
      -- CP-element group 226: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_Update/req
      -- 
    ack_2630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1126_inst_ack_0, ack => zeropad_CP_920_elements(226)); -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(226), ack => WPIPE_Zeropad_output_pipe_1126_inst_req_1); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1126_Update/ack
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1126_inst_ack_1, ack => zeropad_CP_920_elements(227)); -- 
    -- CP-element group 228:  join  transition  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	208 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_Sample/req
      -- 
    req_2643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(228), ack => WPIPE_Zeropad_output_pipe_1129_inst_req_0); -- 
    zeropad_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(208) & zeropad_CP_920_elements(227);
      gj_zeropad_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (6) 
      -- CP-element group 229: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_sample_completed_
      -- CP-element group 229: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_update_start_
      -- CP-element group 229: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_Sample/ack
      -- CP-element group 229: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_Update/req
      -- 
    ack_2644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1129_inst_ack_0, ack => zeropad_CP_920_elements(229)); -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(229), ack => WPIPE_Zeropad_output_pipe_1129_inst_req_1); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1129_Update/ack
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1129_inst_ack_1, ack => zeropad_CP_920_elements(230)); -- 
    -- CP-element group 231:  join  transition  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	206 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_Sample/req
      -- 
    req_2657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(231), ack => WPIPE_Zeropad_output_pipe_1132_inst_req_0); -- 
    zeropad_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(206) & zeropad_CP_920_elements(230);
      gj_zeropad_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_update_start_
      -- CP-element group 232: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_Sample/ack
      -- CP-element group 232: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_Update/$entry
      -- CP-element group 232: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_Update/req
      -- 
    ack_2658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1132_inst_ack_0, ack => zeropad_CP_920_elements(232)); -- 
    req_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(232), ack => WPIPE_Zeropad_output_pipe_1132_inst_req_1); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1132_Update/ack
      -- 
    ack_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1132_inst_ack_1, ack => zeropad_CP_920_elements(233)); -- 
    -- CP-element group 234:  join  transition  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	204 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_Sample/req
      -- 
    req_2671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(234), ack => WPIPE_Zeropad_output_pipe_1135_inst_req_0); -- 
    zeropad_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(204) & zeropad_CP_920_elements(233);
      gj_zeropad_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_update_start_
      -- CP-element group 235: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_Update/req
      -- 
    ack_2672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1135_inst_ack_0, ack => zeropad_CP_920_elements(235)); -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(235), ack => WPIPE_Zeropad_output_pipe_1135_inst_req_1); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1135_Update/ack
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1135_inst_ack_1, ack => zeropad_CP_920_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	202 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_Sample/req
      -- 
    req_2685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(237), ack => WPIPE_Zeropad_output_pipe_1138_inst_req_0); -- 
    zeropad_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(202) & zeropad_CP_920_elements(236);
      gj_zeropad_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_sample_completed_
      -- CP-element group 238: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_update_start_
      -- CP-element group 238: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_Sample/ack
      -- CP-element group 238: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_Update/req
      -- 
    ack_2686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1138_inst_ack_0, ack => zeropad_CP_920_elements(238)); -- 
    req_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(238), ack => WPIPE_Zeropad_output_pipe_1138_inst_req_1); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/WPIPE_Zeropad_output_pipe_1138_Update/ack
      -- 
    ack_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1138_inst_ack_1, ack => zeropad_CP_920_elements(239)); -- 
    -- CP-element group 240:  branch  join  transition  place  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	195 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (10) 
      -- CP-element group 240: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151__exit__
      -- CP-element group 240: 	 branch_block_stmt_316/if_stmt_1152__entry__
      -- CP-element group 240: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/$exit
      -- CP-element group 240: 	 branch_block_stmt_316/if_stmt_1152_dead_link/$entry
      -- CP-element group 240: 	 branch_block_stmt_316/if_stmt_1152_eval_test/$entry
      -- CP-element group 240: 	 branch_block_stmt_316/if_stmt_1152_eval_test/$exit
      -- CP-element group 240: 	 branch_block_stmt_316/if_stmt_1152_eval_test/branch_req
      -- CP-element group 240: 	 branch_block_stmt_316/R_exitcond8_1153_place
      -- CP-element group 240: 	 branch_block_stmt_316/if_stmt_1152_if_link/$entry
      -- CP-element group 240: 	 branch_block_stmt_316/if_stmt_1152_else_link/$entry
      -- 
    branch_req_2699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(240), ack => if_stmt_1152_branch_req_0); -- 
    zeropad_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(195) & zeropad_CP_920_elements(239);
      gj_zeropad_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  merge  transition  place  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	263 
    -- CP-element group 241:  members (13) 
      -- CP-element group 241: 	 branch_block_stmt_316/merge_stmt_1158_PhiReqMerge
      -- CP-element group 241: 	 branch_block_stmt_316/merge_stmt_1158__exit__
      -- CP-element group 241: 	 branch_block_stmt_316/forx_xend287x_xloopexit_forx_xend287
      -- CP-element group 241: 	 branch_block_stmt_316/forx_xbody215_forx_xend287x_xloopexit_PhiReq/$entry
      -- CP-element group 241: 	 branch_block_stmt_316/forx_xbody215_forx_xend287x_xloopexit_PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_316/merge_stmt_1158_PhiAck/$entry
      -- CP-element group 241: 	 branch_block_stmt_316/merge_stmt_1158_PhiAck/$exit
      -- CP-element group 241: 	 branch_block_stmt_316/merge_stmt_1158_PhiAck/dummy
      -- CP-element group 241: 	 branch_block_stmt_316/forx_xend287x_xloopexit_forx_xend287_PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_316/forx_xend287x_xloopexit_forx_xend287_PhiReq/$entry
      -- CP-element group 241: 	 branch_block_stmt_316/if_stmt_1152_if_link/$exit
      -- CP-element group 241: 	 branch_block_stmt_316/if_stmt_1152_if_link/if_choice_transition
      -- CP-element group 241: 	 branch_block_stmt_316/forx_xbody215_forx_xend287x_xloopexit
      -- 
    if_choice_transition_2704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1152_branch_ack_1, ack => zeropad_CP_920_elements(241)); -- 
    -- CP-element group 242:  fork  transition  place  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	258 
    -- CP-element group 242: 	259 
    -- CP-element group 242:  members (12) 
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/$entry
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/$entry
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/$entry
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/$entry
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/Sample/rr
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/Update/cr
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/$entry
      -- CP-element group 242: 	 branch_block_stmt_316/if_stmt_1152_else_link/$exit
      -- CP-element group 242: 	 branch_block_stmt_316/if_stmt_1152_else_link/else_choice_transition
      -- CP-element group 242: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215
      -- 
    else_choice_transition_2708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1152_branch_ack_0, ack => zeropad_CP_920_elements(242)); -- 
    rr_2906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(242), ack => type_cast_1028_inst_req_0); -- 
    cr_2911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(242), ack => type_cast_1028_inst_req_1); -- 
    -- CP-element group 243:  merge  branch  transition  place  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	119 
    -- CP-element group 243: 	69 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	70 
    -- CP-element group 243: 	71 
    -- CP-element group 243:  members (17) 
      -- CP-element group 243: 	 branch_block_stmt_316/merge_stmt_525__exit__
      -- CP-element group 243: 	 branch_block_stmt_316/assign_stmt_531__entry__
      -- CP-element group 243: 	 branch_block_stmt_316/assign_stmt_531__exit__
      -- CP-element group 243: 	 branch_block_stmt_316/if_stmt_532__entry__
      -- CP-element group 243: 	 branch_block_stmt_316/assign_stmt_531/$entry
      -- CP-element group 243: 	 branch_block_stmt_316/assign_stmt_531/$exit
      -- CP-element group 243: 	 branch_block_stmt_316/if_stmt_532_dead_link/$entry
      -- CP-element group 243: 	 branch_block_stmt_316/if_stmt_532_eval_test/$entry
      -- CP-element group 243: 	 branch_block_stmt_316/if_stmt_532_eval_test/$exit
      -- CP-element group 243: 	 branch_block_stmt_316/if_stmt_532_eval_test/branch_req
      -- CP-element group 243: 	 branch_block_stmt_316/R_cmp123292_533_place
      -- CP-element group 243: 	 branch_block_stmt_316/if_stmt_532_if_link/$entry
      -- CP-element group 243: 	 branch_block_stmt_316/if_stmt_532_else_link/$entry
      -- CP-element group 243: 	 branch_block_stmt_316/merge_stmt_525_PhiReqMerge
      -- CP-element group 243: 	 branch_block_stmt_316/merge_stmt_525_PhiAck/$entry
      -- CP-element group 243: 	 branch_block_stmt_316/merge_stmt_525_PhiAck/$exit
      -- CP-element group 243: 	 branch_block_stmt_316/merge_stmt_525_PhiAck/dummy
      -- 
    branch_req_1440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(243), ack => if_stmt_532_branch_req_0); -- 
    zeropad_CP_920_elements(243) <= OrReduce(zeropad_CP_920_elements(119) & zeropad_CP_920_elements(69));
    -- CP-element group 244:  transition  output  delay-element  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	78 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	248 
    -- CP-element group 244:  members (5) 
      -- CP-element group 244: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/$exit
      -- CP-element group 244: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_586_konst_delay_trans
      -- CP-element group 244: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_req
      -- CP-element group 244: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody_PhiReq/phi_stmt_582/$exit
      -- CP-element group 244: 	 branch_block_stmt_316/bbx_xnph298_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_582_req_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_582_req_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(244), ack => phi_stmt_582_req_0); -- 
    -- Element group zeropad_CP_920_elements(244) is a control-delay.
    cp_element_244_delay: control_delay_element  generic map(name => " 244_delay", delay_value => 1)  port map(req => zeropad_CP_920_elements(78), ack => zeropad_CP_920_elements(244), clk => clk, reset =>reset);
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	120 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (2) 
      -- CP-element group 245: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/Sample/ra
      -- CP-element group 245: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/Sample/$exit
      -- 
    ra_2776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_588_inst_ack_0, ack => zeropad_CP_920_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	120 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/Update/ca
      -- CP-element group 246: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/Update/$exit
      -- 
    ca_2781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_588_inst_ack_1, ack => zeropad_CP_920_elements(246)); -- 
    -- CP-element group 247:  join  transition  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 247: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/$exit
      -- CP-element group 247: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_req
      -- CP-element group 247: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/SplitProtocol/$exit
      -- CP-element group 247: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/type_cast_588/$exit
      -- CP-element group 247: 	 branch_block_stmt_316/forx_xbody_forx_xbody_PhiReq/phi_stmt_582/phi_stmt_582_sources/$exit
      -- 
    phi_stmt_582_req_2782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_582_req_2782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(247), ack => phi_stmt_582_req_1); -- 
    zeropad_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(245) & zeropad_CP_920_elements(246);
      gj_zeropad_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  merge  transition  place  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	244 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (2) 
      -- CP-element group 248: 	 branch_block_stmt_316/merge_stmt_581_PhiAck/$entry
      -- CP-element group 248: 	 branch_block_stmt_316/merge_stmt_581_PhiReqMerge
      -- 
    zeropad_CP_920_elements(248) <= OrReduce(zeropad_CP_920_elements(244) & zeropad_CP_920_elements(247));
    -- CP-element group 249:  fork  transition  place  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	86 
    -- CP-element group 249: 	94 
    -- CP-element group 249: 	83 
    -- CP-element group 249: 	82 
    -- CP-element group 249: 	79 
    -- CP-element group 249: 	80 
    -- CP-element group 249: 	90 
    -- CP-element group 249: 	117 
    -- CP-element group 249: 	114 
    -- CP-element group 249: 	106 
    -- CP-element group 249: 	110 
    -- CP-element group 249: 	98 
    -- CP-element group 249: 	102 
    -- CP-element group 249:  members (56) 
      -- CP-element group 249: 	 branch_block_stmt_316/merge_stmt_581__exit__
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746__entry__
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_resized_2
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_scaled_2
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_computed_2
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_resize_2/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_resize_2/$exit
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_resize_2/index_resize_req
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_resize_2/index_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_scale_2/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_scale_2/$exit
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_scale_2/scale_rename_req
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_index_scale_2/scale_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_update_start
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_Sample/req
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/array_obj_ref_596_final_index_sum_regn_Update/req
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/addr_of_597_complete/req
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/RPIPE_Zeropad_input_pipe_600_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_604_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_617_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_635_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_653_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_671_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_689_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_707_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/type_cast_725_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_update_start_
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Update/word_access_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Update/word_access_complete/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_316/assign_stmt_598_to_assign_stmt_746/ptr_deref_733_Update/word_access_complete/word_0/cr
      -- CP-element group 249: 	 branch_block_stmt_316/merge_stmt_581_PhiAck/phi_stmt_582_ack
      -- CP-element group 249: 	 branch_block_stmt_316/merge_stmt_581_PhiAck/$exit
      -- 
    phi_stmt_582_ack_2787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_582_ack_0, ack => zeropad_CP_920_elements(249)); -- 
    req_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => array_obj_ref_596_index_offset_req_0); -- 
    req_1529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => array_obj_ref_596_index_offset_req_1); -- 
    req_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => addr_of_597_final_reg_req_1); -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => RPIPE_Zeropad_input_pipe_600_inst_req_0); -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => type_cast_604_inst_req_1); -- 
    cr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => type_cast_617_inst_req_1); -- 
    cr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => type_cast_635_inst_req_1); -- 
    cr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => type_cast_653_inst_req_1); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => type_cast_671_inst_req_1); -- 
    cr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => type_cast_689_inst_req_1); -- 
    cr_1740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => type_cast_707_inst_req_1); -- 
    cr_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => type_cast_725_inst_req_1); -- 
    cr_1818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(249), ack => ptr_deref_733_store_0_req_1); -- 
    -- CP-element group 250:  transition  output  delay-element  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	127 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	254 
    -- CP-element group 250:  members (5) 
      -- CP-element group 250: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_req
      -- CP-element group 250: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801_konst_delay_trans
      -- CP-element group 250: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/$exit
      -- CP-element group 250: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125_PhiReq/phi_stmt_797/$exit
      -- CP-element group 250: 	 branch_block_stmt_316/bbx_xnph294_forx_xbody125_PhiReq/$exit
      -- 
    phi_stmt_797_req_2810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_797_req_2810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(250), ack => phi_stmt_797_req_0); -- 
    -- Element group zeropad_CP_920_elements(250) is a control-delay.
    cp_element_250_delay: control_delay_element  generic map(name => " 250_delay", delay_value => 1)  port map(req => zeropad_CP_920_elements(127), ack => zeropad_CP_920_elements(250), clk => clk, reset =>reset);
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	136 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/Sample/ra
      -- 
    ra_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_803_inst_ack_0, ack => zeropad_CP_920_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	136 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (2) 
      -- CP-element group 252: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/Update/ca
      -- 
    ca_2835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_803_inst_ack_1, ack => zeropad_CP_920_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/$exit
      -- CP-element group 253: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/$exit
      -- CP-element group 253: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/$exit
      -- CP-element group 253: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/$exit
      -- CP-element group 253: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_803/SplitProtocol/$exit
      -- CP-element group 253: 	 branch_block_stmt_316/forx_xbody125_forx_xbody125_PhiReq/phi_stmt_797/phi_stmt_797_req
      -- 
    phi_stmt_797_req_2836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_797_req_2836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(253), ack => phi_stmt_797_req_1); -- 
    zeropad_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(251) & zeropad_CP_920_elements(252);
      gj_zeropad_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  merge  transition  place  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	250 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_316/merge_stmt_796_PhiReqMerge
      -- CP-element group 254: 	 branch_block_stmt_316/merge_stmt_796_PhiAck/$entry
      -- 
    zeropad_CP_920_elements(254) <= OrReduce(zeropad_CP_920_elements(250) & zeropad_CP_920_elements(253));
    -- CP-element group 255:  fork  transition  place  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	131 
    -- CP-element group 255: 	128 
    -- CP-element group 255: 	129 
    -- CP-element group 255: 	133 
    -- CP-element group 255:  members (29) 
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_update_start_
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_complete/req
      -- CP-element group 255: 	 branch_block_stmt_316/merge_stmt_796__exit__
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829__entry__
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Update/word_access_complete/word_0/cr
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_complete/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Update/word_access_complete/word_0/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Update/word_access_complete/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/ptr_deref_815_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/addr_of_812_update_start_
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_resized_2
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_scaled_2
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_computed_2
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_resize_2/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_resize_2/$exit
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_resize_2/index_resize_req
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_resize_2/index_resize_ack
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_scale_2/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_scale_2/$exit
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_scale_2/scale_rename_req
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_index_scale_2/scale_rename_ack
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_update_start
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_Sample/req
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_316/assign_stmt_813_to_assign_stmt_829/array_obj_ref_811_final_index_sum_regn_Update/req
      -- CP-element group 255: 	 branch_block_stmt_316/merge_stmt_796_PhiAck/phi_stmt_797_ack
      -- CP-element group 255: 	 branch_block_stmt_316/merge_stmt_796_PhiAck/$exit
      -- 
    phi_stmt_797_ack_2841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_797_ack_0, ack => zeropad_CP_920_elements(255)); -- 
    req_1931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(255), ack => addr_of_812_final_reg_req_1); -- 
    cr_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(255), ack => ptr_deref_815_store_0_req_1); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(255), ack => array_obj_ref_811_index_offset_req_0); -- 
    req_1916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(255), ack => array_obj_ref_811_index_offset_req_1); -- 
    -- CP-element group 256:  merge  fork  transition  place  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	71 
    -- CP-element group 256: 	135 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	140 
    -- CP-element group 256: 	137 
    -- CP-element group 256: 	138 
    -- CP-element group 256:  members (16) 
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/$entry
      -- CP-element group 256: 	 branch_block_stmt_316/merge_stmt_838_PhiReqMerge
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_update_start_
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_Sample/crr
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/call_stmt_841_Update/ccr
      -- CP-element group 256: 	 branch_block_stmt_316/merge_stmt_838__exit__
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847__entry__
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_update_start_
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_Update/cr
      -- CP-element group 256: 	 branch_block_stmt_316/call_stmt_841_to_assign_stmt_847/type_cast_846_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_316/merge_stmt_838_PhiAck/dummy
      -- CP-element group 256: 	 branch_block_stmt_316/merge_stmt_838_PhiAck/$exit
      -- CP-element group 256: 	 branch_block_stmt_316/merge_stmt_838_PhiAck/$entry
      -- 
    crr_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(256), ack => call_stmt_841_call_req_0); -- 
    ccr_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(256), ack => call_stmt_841_call_req_1); -- 
    cr_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(256), ack => type_cast_846_inst_req_1); -- 
    zeropad_CP_920_elements(256) <= OrReduce(zeropad_CP_920_elements(71) & zeropad_CP_920_elements(135));
    -- CP-element group 257:  transition  output  delay-element  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	194 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	261 
    -- CP-element group 257:  members (5) 
      -- CP-element group 257: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_req
      -- CP-element group 257: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1026_konst_delay_trans
      -- CP-element group 257: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/$exit
      -- CP-element group 257: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215_PhiReq/phi_stmt_1022/$exit
      -- CP-element group 257: 	 branch_block_stmt_316/bbx_xnph_forx_xbody215_PhiReq/$exit
      -- 
    phi_stmt_1022_req_2887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1022_req_2887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(257), ack => phi_stmt_1022_req_0); -- 
    -- Element group zeropad_CP_920_elements(257) is a control-delay.
    cp_element_257_delay: control_delay_element  generic map(name => " 257_delay", delay_value => 1)  port map(req => zeropad_CP_920_elements(194), ack => zeropad_CP_920_elements(257), clk => clk, reset =>reset);
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	242 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/Sample/ra
      -- 
    ra_2907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1028_inst_ack_0, ack => zeropad_CP_920_elements(258)); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	242 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (2) 
      -- CP-element group 259: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/Update/ca
      -- 
    ca_2912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1028_inst_ack_1, ack => zeropad_CP_920_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/$exit
      -- CP-element group 260: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/$exit
      -- CP-element group 260: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/$exit
      -- CP-element group 260: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/$exit
      -- CP-element group 260: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_sources/type_cast_1028/SplitProtocol/$exit
      -- CP-element group 260: 	 branch_block_stmt_316/forx_xbody215_forx_xbody215_PhiReq/phi_stmt_1022/phi_stmt_1022_req
      -- 
    phi_stmt_1022_req_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1022_req_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(260), ack => phi_stmt_1022_req_1); -- 
    zeropad_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_920_elements(258) & zeropad_CP_920_elements(259);
      gj_zeropad_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_920_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  merge  transition  place  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	257 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (2) 
      -- CP-element group 261: 	 branch_block_stmt_316/merge_stmt_1021_PhiReqMerge
      -- CP-element group 261: 	 branch_block_stmt_316/merge_stmt_1021_PhiAck/$entry
      -- 
    zeropad_CP_920_elements(261) <= OrReduce(zeropad_CP_920_elements(257) & zeropad_CP_920_elements(260));
    -- CP-element group 262:  fork  transition  place  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	195 
    -- CP-element group 262: 	196 
    -- CP-element group 262: 	198 
    -- CP-element group 262: 	200 
    -- CP-element group 262: 	202 
    -- CP-element group 262: 	204 
    -- CP-element group 262: 	206 
    -- CP-element group 262: 	208 
    -- CP-element group 262: 	210 
    -- CP-element group 262: 	212 
    -- CP-element group 262: 	214 
    -- CP-element group 262: 	216 
    -- CP-element group 262:  members (53) 
      -- CP-element group 262: 	 branch_block_stmt_316/merge_stmt_1021__exit__
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151__entry__
      -- CP-element group 262: 	 branch_block_stmt_316/merge_stmt_1021_PhiAck/$exit
      -- CP-element group 262: 	 branch_block_stmt_316/merge_stmt_1021_PhiAck/phi_stmt_1022_ack
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_resized_2
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_scaled_2
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_computed_2
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_resize_2/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_resize_2/$exit
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_resize_2/index_resize_req
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_resize_2/index_resize_ack
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_scale_2/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_scale_2/$exit
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_scale_2/scale_rename_req
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_index_scale_2/scale_rename_ack
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_update_start
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_Sample/req
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/array_obj_ref_1036_final_index_sum_regn_Update/req
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_complete/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/addr_of_1037_complete/req
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/word_access_complete/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/word_access_complete/word_0/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/ptr_deref_1041_Update/word_access_complete/word_0/cr
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1045_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1055_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1065_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1075_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1085_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1095_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1105_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_update_start_
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_316/assign_stmt_1038_to_assign_stmt_1151/type_cast_1115_Update/cr
      -- 
    phi_stmt_1022_ack_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1022_ack_0, ack => zeropad_CP_920_elements(262)); -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => array_obj_ref_1036_index_offset_req_0); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => array_obj_ref_1036_index_offset_req_1); -- 
    req_2416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => addr_of_1037_final_reg_req_1); -- 
    cr_2461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => ptr_deref_1041_load_0_req_1); -- 
    cr_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => type_cast_1045_inst_req_1); -- 
    cr_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => type_cast_1055_inst_req_1); -- 
    cr_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => type_cast_1065_inst_req_1); -- 
    cr_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => type_cast_1075_inst_req_1); -- 
    cr_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => type_cast_1085_inst_req_1); -- 
    cr_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => type_cast_1095_inst_req_1); -- 
    cr_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => type_cast_1105_inst_req_1); -- 
    cr_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_920_elements(262), ack => type_cast_1115_inst_req_1); -- 
    -- CP-element group 263:  merge  transition  place  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	187 
    -- CP-element group 263: 	241 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (16) 
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1162_PhiReqMerge
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1160_PhiReqMerge
      -- CP-element group 263: 	 $exit
      -- CP-element group 263: 	 branch_block_stmt_316/$exit
      -- CP-element group 263: 	 branch_block_stmt_316/branch_block_stmt_316__exit__
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1160__exit__
      -- CP-element group 263: 	 branch_block_stmt_316/return__
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1162__exit__
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1162_PhiAck/dummy
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1162_PhiAck/$exit
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1162_PhiAck/$entry
      -- CP-element group 263: 	 branch_block_stmt_316/return___PhiReq/$exit
      -- CP-element group 263: 	 branch_block_stmt_316/return___PhiReq/$entry
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1160_PhiAck/dummy
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1160_PhiAck/$exit
      -- CP-element group 263: 	 branch_block_stmt_316/merge_stmt_1160_PhiAck/$entry
      -- 
    zeropad_CP_920_elements(263) <= OrReduce(zeropad_CP_920_elements(187) & zeropad_CP_920_elements(241));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_ix_x0297_595_resized : std_logic_vector(14 downto 0);
    signal R_ix_x0297_595_scaled : std_logic_vector(14 downto 0);
    signal R_ix_x1293_810_resized : std_logic_vector(14 downto 0);
    signal R_ix_x1293_810_scaled : std_logic_vector(14 downto 0);
    signal R_ix_x2290_1035_resized : std_logic_vector(14 downto 0);
    signal R_ix_x2290_1035_scaled : std_logic_vector(14 downto 0);
    signal add103_695 : std_logic_vector(63 downto 0);
    signal add109_713 : std_logic_vector(63 downto 0);
    signal add115_731 : std_logic_vector(63 downto 0);
    signal add12_366 : std_logic_vector(15 downto 0);
    signal add21_391 : std_logic_vector(15 downto 0);
    signal add30_416 : std_logic_vector(15 downto 0);
    signal add39_441 : std_logic_vector(15 downto 0);
    signal add48_466 : std_logic_vector(15 downto 0);
    signal add79_623 : std_logic_vector(63 downto 0);
    signal add85_641 : std_logic_vector(63 downto 0);
    signal add91_659 : std_logic_vector(63 downto 0);
    signal add97_677 : std_logic_vector(63 downto 0);
    signal add_341 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1036_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_1036_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_1036_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1036_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1036_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1036_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_1036_root_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_596_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_596_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_596_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_596_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_596_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_596_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_596_root_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_811_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_811_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_811_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_811_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_811_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_811_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_811_root_address : std_logic_vector(14 downto 0);
    signal arrayidx127_813 : std_logic_vector(31 downto 0);
    signal arrayidx219_1038 : std_logic_vector(31 downto 0);
    signal arrayidx_598 : std_logic_vector(31 downto 0);
    signal call100_686 : std_logic_vector(7 downto 0);
    signal call106_704 : std_logic_vector(7 downto 0);
    signal call10_357 : std_logic_vector(7 downto 0);
    signal call112_722 : std_logic_vector(7 downto 0);
    signal call133_841 : std_logic_vector(63 downto 0);
    signal call142_862 : std_logic_vector(63 downto 0);
    signal call14_369 : std_logic_vector(7 downto 0);
    signal call19_382 : std_logic_vector(7 downto 0);
    signal call23_394 : std_logic_vector(7 downto 0);
    signal call28_407 : std_logic_vector(7 downto 0);
    signal call2_332 : std_logic_vector(7 downto 0);
    signal call32_419 : std_logic_vector(7 downto 0);
    signal call37_432 : std_logic_vector(7 downto 0);
    signal call41_444 : std_logic_vector(7 downto 0);
    signal call46_457 : std_logic_vector(7 downto 0);
    signal call5_344 : std_logic_vector(7 downto 0);
    signal call72_601 : std_logic_vector(7 downto 0);
    signal call76_614 : std_logic_vector(7 downto 0);
    signal call82_632 : std_logic_vector(7 downto 0);
    signal call88_650 : std_logic_vector(7 downto 0);
    signal call94_668 : std_logic_vector(7 downto 0);
    signal call_319 : std_logic_vector(7 downto 0);
    signal cmp123292_531 : std_logic_vector(0 downto 0);
    signal cmp296_516 : std_logic_vector(0 downto 0);
    signal conv102_690 : std_logic_vector(63 downto 0);
    signal conv108_708 : std_logic_vector(63 downto 0);
    signal conv114_726 : std_logic_vector(63 downto 0);
    signal conv11_361 : std_logic_vector(15 downto 0);
    signal conv134_847 : std_logic_vector(63 downto 0);
    signal conv143_867 : std_logic_vector(63 downto 0);
    signal conv149_876 : std_logic_vector(7 downto 0);
    signal conv155_886 : std_logic_vector(7 downto 0);
    signal conv161_896 : std_logic_vector(7 downto 0);
    signal conv167_906 : std_logic_vector(7 downto 0);
    signal conv173_916 : std_logic_vector(7 downto 0);
    signal conv179_926 : std_logic_vector(7 downto 0);
    signal conv17_373 : std_logic_vector(15 downto 0);
    signal conv185_936 : std_logic_vector(7 downto 0);
    signal conv191_946 : std_logic_vector(7 downto 0);
    signal conv1_323 : std_logic_vector(15 downto 0);
    signal conv20_386 : std_logic_vector(15 downto 0);
    signal conv224_1046 : std_logic_vector(7 downto 0);
    signal conv230_1056 : std_logic_vector(7 downto 0);
    signal conv236_1066 : std_logic_vector(7 downto 0);
    signal conv242_1076 : std_logic_vector(7 downto 0);
    signal conv248_1086 : std_logic_vector(7 downto 0);
    signal conv254_1096 : std_logic_vector(7 downto 0);
    signal conv260_1106 : std_logic_vector(7 downto 0);
    signal conv266_1116 : std_logic_vector(7 downto 0);
    signal conv26_398 : std_logic_vector(15 downto 0);
    signal conv29_411 : std_logic_vector(15 downto 0);
    signal conv35_423 : std_logic_vector(15 downto 0);
    signal conv38_436 : std_logic_vector(15 downto 0);
    signal conv3_336 : std_logic_vector(15 downto 0);
    signal conv44_448 : std_logic_vector(15 downto 0);
    signal conv47_461 : std_logic_vector(15 downto 0);
    signal conv53_470 : std_logic_vector(31 downto 0);
    signal conv55_474 : std_logic_vector(31 downto 0);
    signal conv57_478 : std_logic_vector(31 downto 0);
    signal conv61_492 : std_logic_vector(31 downto 0);
    signal conv63_496 : std_logic_vector(31 downto 0);
    signal conv66_500 : std_logic_vector(31 downto 0);
    signal conv73_605 : std_logic_vector(63 downto 0);
    signal conv78_618 : std_logic_vector(63 downto 0);
    signal conv84_636 : std_logic_vector(63 downto 0);
    signal conv8_348 : std_logic_vector(15 downto 0);
    signal conv90_654 : std_logic_vector(63 downto 0);
    signal conv96_672 : std_logic_vector(63 downto 0);
    signal exitcond24_746 : std_logic_vector(0 downto 0);
    signal exitcond8_1151 : std_logic_vector(0 downto 0);
    signal exitcond_829 : std_logic_vector(0 downto 0);
    signal inc130_824 : std_logic_vector(31 downto 0);
    signal inc286_1146 : std_logic_vector(31 downto 0);
    signal inc_741 : std_logic_vector(31 downto 0);
    signal ix_x0297_582 : std_logic_vector(31 downto 0);
    signal ix_x1293_797 : std_logic_vector(31 downto 0);
    signal ix_x2290_1022 : std_logic_vector(31 downto 0);
    signal mul58_488 : std_logic_vector(31 downto 0);
    signal mul64_505 : std_logic_vector(31 downto 0);
    signal mul67_510 : std_logic_vector(31 downto 0);
    signal mul_483 : std_logic_vector(31 downto 0);
    signal ptr_deref_1041_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1041_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_1041_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_1041_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_1041_word_offset_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_733_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_733_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_733_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_733_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_733_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_733_word_offset_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_815_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_815_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_815_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_815_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_815_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_815_word_offset_0 : std_logic_vector(14 downto 0);
    signal shl105_701 : std_logic_vector(63 downto 0);
    signal shl111_719 : std_logic_vector(63 downto 0);
    signal shl18_379 : std_logic_vector(15 downto 0);
    signal shl27_404 : std_logic_vector(15 downto 0);
    signal shl36_429 : std_logic_vector(15 downto 0);
    signal shl45_454 : std_logic_vector(15 downto 0);
    signal shl75_611 : std_logic_vector(63 downto 0);
    signal shl81_629 : std_logic_vector(63 downto 0);
    signal shl87_647 : std_logic_vector(63 downto 0);
    signal shl93_665 : std_logic_vector(63 downto 0);
    signal shl99_683 : std_logic_vector(63 downto 0);
    signal shl9_354 : std_logic_vector(15 downto 0);
    signal shl_329 : std_logic_vector(15 downto 0);
    signal shr152_882 : std_logic_vector(63 downto 0);
    signal shr158_892 : std_logic_vector(63 downto 0);
    signal shr164_902 : std_logic_vector(63 downto 0);
    signal shr170_912 : std_logic_vector(63 downto 0);
    signal shr176_922 : std_logic_vector(63 downto 0);
    signal shr182_932 : std_logic_vector(63 downto 0);
    signal shr188_942 : std_logic_vector(63 downto 0);
    signal shr227_1052 : std_logic_vector(63 downto 0);
    signal shr233_1062 : std_logic_vector(63 downto 0);
    signal shr239_1072 : std_logic_vector(63 downto 0);
    signal shr245_1082 : std_logic_vector(63 downto 0);
    signal shr251_1092 : std_logic_vector(63 downto 0);
    signal shr257_1102 : std_logic_vector(63 downto 0);
    signal shr263_1112 : std_logic_vector(63 downto 0);
    signal sub_872 : std_logic_vector(63 downto 0);
    signal tmp10_761 : std_logic_vector(31 downto 0);
    signal tmp11_766 : std_logic_vector(31 downto 0);
    signal tmp12_770 : std_logic_vector(31 downto 0);
    signal tmp13_775 : std_logic_vector(31 downto 0);
    signal tmp14_781 : std_logic_vector(31 downto 0);
    signal tmp15_787 : std_logic_vector(0 downto 0);
    signal tmp16_542 : std_logic_vector(31 downto 0);
    signal tmp17_546 : std_logic_vector(31 downto 0);
    signal tmp18_551 : std_logic_vector(31 downto 0);
    signal tmp19_555 : std_logic_vector(31 downto 0);
    signal tmp1_986 : std_logic_vector(31 downto 0);
    signal tmp20_560 : std_logic_vector(31 downto 0);
    signal tmp21_566 : std_logic_vector(31 downto 0);
    signal tmp220_1042 : std_logic_vector(63 downto 0);
    signal tmp22_572 : std_logic_vector(0 downto 0);
    signal tmp2_991 : std_logic_vector(31 downto 0);
    signal tmp3_995 : std_logic_vector(31 downto 0);
    signal tmp4_1000 : std_logic_vector(31 downto 0);
    signal tmp5_1006 : std_logic_vector(31 downto 0);
    signal tmp6_1012 : std_logic_vector(0 downto 0);
    signal tmp9_757 : std_logic_vector(31 downto 0);
    signal tmp_982 : std_logic_vector(31 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1010_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1017_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1026_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1028_wire : std_logic_vector(31 downto 0);
    signal type_cast_1050_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1060_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1070_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1080_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1090_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1100_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1110_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_327_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_352_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_377_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_402_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_427_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_452_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_514_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_529_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_564_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_570_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_577_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_586_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_588_wire : std_logic_vector(31 downto 0);
    signal type_cast_609_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_627_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_645_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_663_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_681_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_699_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_717_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_739_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_779_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_785_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_792_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_801_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_803_wire : std_logic_vector(31 downto 0);
    signal type_cast_817_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_822_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_845_wire : std_logic_vector(63 downto 0);
    signal type_cast_856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_858_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_865_wire : std_logic_vector(63 downto 0);
    signal type_cast_880_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_900_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_910_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_930_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_940_wire_constant : std_logic_vector(63 downto 0);
    signal umax23_579 : std_logic_vector(31 downto 0);
    signal umax7_1019 : std_logic_vector(31 downto 0);
    signal umax_794 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1036_constant_part_of_offset <= "100000000000000";
    array_obj_ref_1036_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_1036_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_1036_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_1036_resized_base_address <= "000000000000000";
    array_obj_ref_596_constant_part_of_offset <= "000000000000000";
    array_obj_ref_596_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_596_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_596_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_596_resized_base_address <= "000000000000000";
    array_obj_ref_811_constant_part_of_offset <= "100000000000000";
    array_obj_ref_811_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_811_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_811_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_811_resized_base_address <= "000000000000000";
    ptr_deref_1041_word_offset_0 <= "000000000000000";
    ptr_deref_733_word_offset_0 <= "000000000000000";
    ptr_deref_815_word_offset_0 <= "000000000000000";
    type_cast_1004_wire_constant <= "00000000000000000000000000000011";
    type_cast_1010_wire_constant <= "00000000000000000000000000000001";
    type_cast_1017_wire_constant <= "00000000000000000000000000000001";
    type_cast_1026_wire_constant <= "00000000000000000000000000000000";
    type_cast_1050_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1060_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1070_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1080_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1090_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1100_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1110_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1144_wire_constant <= "00000000000000000000000000000001";
    type_cast_327_wire_constant <= "0000000000001000";
    type_cast_352_wire_constant <= "0000000000001000";
    type_cast_377_wire_constant <= "0000000000001000";
    type_cast_402_wire_constant <= "0000000000001000";
    type_cast_427_wire_constant <= "0000000000001000";
    type_cast_452_wire_constant <= "0000000000001000";
    type_cast_514_wire_constant <= "00000000000000000000000000000111";
    type_cast_529_wire_constant <= "00000000000000000000000000000111";
    type_cast_564_wire_constant <= "00000000000000000000000000000011";
    type_cast_570_wire_constant <= "00000000000000000000000000000001";
    type_cast_577_wire_constant <= "00000000000000000000000000000001";
    type_cast_586_wire_constant <= "00000000000000000000000000000000";
    type_cast_609_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_627_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_645_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_663_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_681_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_699_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_717_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_739_wire_constant <= "00000000000000000000000000000001";
    type_cast_779_wire_constant <= "00000000000000000000000000000011";
    type_cast_785_wire_constant <= "00000000000000000000000000000001";
    type_cast_792_wire_constant <= "00000000000000000000000000000001";
    type_cast_801_wire_constant <= "00000000000000000000000000000000";
    type_cast_817_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_822_wire_constant <= "00000000000000000000000000000001";
    type_cast_856_wire_constant <= "00000000";
    type_cast_858_wire_constant <= "00000001";
    type_cast_880_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_890_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_900_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_910_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_920_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_930_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_940_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    phi_stmt_1022: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1026_wire_constant & type_cast_1028_wire;
      req <= phi_stmt_1022_req_0 & phi_stmt_1022_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1022",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1022_ack_0,
          idata => idata,
          odata => ix_x2290_1022,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1022
    phi_stmt_582: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_586_wire_constant & type_cast_588_wire;
      req <= phi_stmt_582_req_0 & phi_stmt_582_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_582",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_582_ack_0,
          idata => idata,
          odata => ix_x0297_582,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_582
    phi_stmt_797: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_801_wire_constant & type_cast_803_wire;
      req <= phi_stmt_797_req_0 & phi_stmt_797_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_797",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_797_ack_0,
          idata => idata,
          odata => ix_x1293_797,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_797
    -- flow-through select operator MUX_1018_inst
    umax7_1019 <= tmp5_1006 when (tmp6_1012(0) /=  '0') else type_cast_1017_wire_constant;
    -- flow-through select operator MUX_578_inst
    umax23_579 <= tmp21_566 when (tmp22_572(0) /=  '0') else type_cast_577_wire_constant;
    -- flow-through select operator MUX_793_inst
    umax_794 <= tmp14_781 when (tmp15_787(0) /=  '0') else type_cast_792_wire_constant;
    addr_of_1037_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1037_final_reg_req_0;
      addr_of_1037_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1037_final_reg_req_1;
      addr_of_1037_final_reg_ack_1<= rack(0);
      addr_of_1037_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1037_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1036_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx219_1038,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_597_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_597_final_reg_req_0;
      addr_of_597_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_597_final_reg_req_1;
      addr_of_597_final_reg_ack_1<= rack(0);
      addr_of_597_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_597_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_596_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_812_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_812_final_reg_req_0;
      addr_of_812_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_812_final_reg_req_1;
      addr_of_812_final_reg_ack_1<= rack(0);
      addr_of_812_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_812_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_811_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx127_813,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1028_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1028_inst_req_0;
      type_cast_1028_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1028_inst_req_1;
      type_cast_1028_inst_ack_1<= rack(0);
      type_cast_1028_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1028_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc286_1146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1028_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1045_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1045_inst_req_0;
      type_cast_1045_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1045_inst_req_1;
      type_cast_1045_inst_ack_1<= rack(0);
      type_cast_1045_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1045_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp220_1042,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv224_1046,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1055_inst_req_0;
      type_cast_1055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1055_inst_req_1;
      type_cast_1055_inst_ack_1<= rack(0);
      type_cast_1055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr227_1052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_1056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1065_inst_req_0;
      type_cast_1065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1065_inst_req_1;
      type_cast_1065_inst_ack_1<= rack(0);
      type_cast_1065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr233_1062,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv236_1066,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1075_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1075_inst_req_0;
      type_cast_1075_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1075_inst_req_1;
      type_cast_1075_inst_ack_1<= rack(0);
      type_cast_1075_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1075_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr239_1072,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv242_1076,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1085_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1085_inst_req_0;
      type_cast_1085_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1085_inst_req_1;
      type_cast_1085_inst_ack_1<= rack(0);
      type_cast_1085_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1085_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr245_1082,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv248_1086,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1095_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1095_inst_req_0;
      type_cast_1095_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1095_inst_req_1;
      type_cast_1095_inst_ack_1<= rack(0);
      type_cast_1095_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1095_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr251_1092,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv254_1096,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1105_inst_req_0;
      type_cast_1105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1105_inst_req_1;
      type_cast_1105_inst_ack_1<= rack(0);
      type_cast_1105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr257_1102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv260_1106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1115_inst_req_0;
      type_cast_1115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1115_inst_req_1;
      type_cast_1115_inst_ack_1<= rack(0);
      type_cast_1115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr263_1112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv266_1116,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_322_inst_req_0;
      type_cast_322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_322_inst_req_1;
      type_cast_322_inst_ack_1<= rack(0);
      type_cast_322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_323,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_335_inst_req_0;
      type_cast_335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_335_inst_req_1;
      type_cast_335_inst_ack_1<= rack(0);
      type_cast_335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_335_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_347_inst_req_0;
      type_cast_347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_347_inst_req_1;
      type_cast_347_inst_ack_1<= rack(0);
      type_cast_347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_344,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_348,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_360_inst_req_0;
      type_cast_360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_360_inst_req_1;
      type_cast_360_inst_ack_1<= rack(0);
      type_cast_360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_372_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_372_inst_req_0;
      type_cast_372_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_372_inst_req_1;
      type_cast_372_inst_ack_1<= rack(0);
      type_cast_372_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_372_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_369,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_373,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_385_inst_req_0;
      type_cast_385_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_385_inst_req_1;
      type_cast_385_inst_ack_1<= rack(0);
      type_cast_385_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_385_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_397_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_397_inst_req_0;
      type_cast_397_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_397_inst_req_1;
      type_cast_397_inst_ack_1<= rack(0);
      type_cast_397_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_397_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_394,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_398,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_410_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_410_inst_req_0;
      type_cast_410_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_410_inst_req_1;
      type_cast_410_inst_ack_1<= rack(0);
      type_cast_410_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_410_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_407,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_411,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_422_inst_req_0;
      type_cast_422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_422_inst_req_1;
      type_cast_422_inst_ack_1<= rack(0);
      type_cast_422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_423,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_435_inst_req_0;
      type_cast_435_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_435_inst_req_1;
      type_cast_435_inst_ack_1<= rack(0);
      type_cast_435_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_435_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_432,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_447_inst_req_0;
      type_cast_447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_447_inst_req_1;
      type_cast_447_inst_ack_1<= rack(0);
      type_cast_447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_447_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_448,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_460_inst_req_0;
      type_cast_460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_460_inst_req_1;
      type_cast_460_inst_ack_1<= rack(0);
      type_cast_460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_461,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_469_inst_req_0;
      type_cast_469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_469_inst_req_1;
      type_cast_469_inst_ack_1<= rack(0);
      type_cast_469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_473_inst_req_0;
      type_cast_473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_473_inst_req_1;
      type_cast_473_inst_ack_1<= rack(0);
      type_cast_473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv55_474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_477_inst_req_0;
      type_cast_477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_477_inst_req_1;
      type_cast_477_inst_ack_1<= rack(0);
      type_cast_477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv57_478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_491_inst_req_0;
      type_cast_491_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_491_inst_req_1;
      type_cast_491_inst_ack_1<= rack(0);
      type_cast_491_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_491_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_492,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_495_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_495_inst_req_0;
      type_cast_495_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_495_inst_req_1;
      type_cast_495_inst_ack_1<= rack(0);
      type_cast_495_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_495_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_496,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_499_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_499_inst_req_0;
      type_cast_499_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_499_inst_req_1;
      type_cast_499_inst_ack_1<= rack(0);
      type_cast_499_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_499_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_500,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_541_inst_req_0;
      type_cast_541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_541_inst_req_1;
      type_cast_541_inst_ack_1<= rack(0);
      type_cast_541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp16_542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_545_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_545_inst_req_0;
      type_cast_545_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_545_inst_req_1;
      type_cast_545_inst_ack_1<= rack(0);
      type_cast_545_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_545_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp17_546,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_554_inst_req_0;
      type_cast_554_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_554_inst_req_1;
      type_cast_554_inst_ack_1<= rack(0);
      type_cast_554_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp19_555,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_588_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_588_inst_req_0;
      type_cast_588_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_588_inst_req_1;
      type_cast_588_inst_ack_1<= rack(0);
      type_cast_588_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_588_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_741,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_588_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_604_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_604_inst_req_0;
      type_cast_604_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_604_inst_req_1;
      type_cast_604_inst_ack_1<= rack(0);
      type_cast_604_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_604_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call72_601,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_605,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_617_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_617_inst_req_0;
      type_cast_617_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_617_inst_req_1;
      type_cast_617_inst_ack_1<= rack(0);
      type_cast_617_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_617_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call76_614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_618,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_635_inst_req_0;
      type_cast_635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_635_inst_req_1;
      type_cast_635_inst_ack_1<= rack(0);
      type_cast_635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_635_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call82_632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_653_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_653_inst_req_0;
      type_cast_653_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_653_inst_req_1;
      type_cast_653_inst_ack_1<= rack(0);
      type_cast_653_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_653_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_650,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_654,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_671_inst_req_0;
      type_cast_671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_671_inst_req_1;
      type_cast_671_inst_ack_1<= rack(0);
      type_cast_671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call94_668,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_689_inst_req_0;
      type_cast_689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_689_inst_req_1;
      type_cast_689_inst_ack_1<= rack(0);
      type_cast_689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call100_686,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv102_690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_707_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_707_inst_req_0;
      type_cast_707_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_707_inst_req_1;
      type_cast_707_inst_ack_1<= rack(0);
      type_cast_707_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_707_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_704,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv108_708,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_725_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_725_inst_req_0;
      type_cast_725_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_725_inst_req_1;
      type_cast_725_inst_ack_1<= rack(0);
      type_cast_725_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_725_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call112_722,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv114_726,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_756_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_756_inst_req_0;
      type_cast_756_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_756_inst_req_1;
      type_cast_756_inst_ack_1<= rack(0);
      type_cast_756_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_756_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp9_757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_760_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_760_inst_req_0;
      type_cast_760_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_760_inst_req_1;
      type_cast_760_inst_ack_1<= rack(0);
      type_cast_760_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_760_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10_761,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_769_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_769_inst_req_0;
      type_cast_769_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_769_inst_req_1;
      type_cast_769_inst_ack_1<= rack(0);
      type_cast_769_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_769_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_770,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_803_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_803_inst_req_0;
      type_cast_803_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_803_inst_req_1;
      type_cast_803_inst_ack_1<= rack(0);
      type_cast_803_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_803_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc130_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_803_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_846_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_846_inst_req_0;
      type_cast_846_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_846_inst_req_1;
      type_cast_846_inst_ack_1<= rack(0);
      type_cast_846_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_846_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_845_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_847,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_866_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_866_inst_req_0;
      type_cast_866_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_866_inst_req_1;
      type_cast_866_inst_ack_1<= rack(0);
      type_cast_866_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_866_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_865_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_867,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_875_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_875_inst_req_0;
      type_cast_875_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_875_inst_req_1;
      type_cast_875_inst_ack_1<= rack(0);
      type_cast_875_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_875_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_876,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_885_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_885_inst_req_0;
      type_cast_885_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_885_inst_req_1;
      type_cast_885_inst_ack_1<= rack(0);
      type_cast_885_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_885_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr152_882,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_886,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_895_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_895_inst_req_0;
      type_cast_895_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_895_inst_req_1;
      type_cast_895_inst_ack_1<= rack(0);
      type_cast_895_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_895_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr158_892,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_896,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_905_inst_req_0;
      type_cast_905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_905_inst_req_1;
      type_cast_905_inst_ack_1<= rack(0);
      type_cast_905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr164_902,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_906,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_915_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_915_inst_req_0;
      type_cast_915_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_915_inst_req_1;
      type_cast_915_inst_ack_1<= rack(0);
      type_cast_915_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_915_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr170_912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_916,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_925_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_925_inst_req_0;
      type_cast_925_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_925_inst_req_1;
      type_cast_925_inst_ack_1<= rack(0);
      type_cast_925_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_925_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr176_922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_926,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_935_inst_req_0;
      type_cast_935_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_935_inst_req_1;
      type_cast_935_inst_ack_1<= rack(0);
      type_cast_935_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_935_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr182_932,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_936,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_945_inst_req_0;
      type_cast_945_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_945_inst_req_1;
      type_cast_945_inst_ack_1<= rack(0);
      type_cast_945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr188_942,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_946,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_981_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_981_inst_req_0;
      type_cast_981_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_981_inst_req_1;
      type_cast_981_inst_ack_1<= rack(0);
      type_cast_981_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_981_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_982,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_985_inst_req_0;
      type_cast_985_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_985_inst_req_1;
      type_cast_985_inst_ack_1<= rack(0);
      type_cast_985_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_986,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_994_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_994_inst_req_0;
      type_cast_994_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_994_inst_req_1;
      type_cast_994_inst_ack_1<= rack(0);
      type_cast_994_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_994_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_995,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1036_index_2_rename
    process(R_ix_x2290_1035_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x2290_1035_resized;
      ov(14 downto 0) := iv;
      R_ix_x2290_1035_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1036_index_2_resize
    process(ix_x2290_1022) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x2290_1022;
      ov := iv(14 downto 0);
      R_ix_x2290_1035_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1036_root_address_inst
    process(array_obj_ref_1036_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1036_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_1036_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_596_index_2_rename
    process(R_ix_x0297_595_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0297_595_resized;
      ov(14 downto 0) := iv;
      R_ix_x0297_595_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_596_index_2_resize
    process(ix_x0297_582) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0297_582;
      ov := iv(14 downto 0);
      R_ix_x0297_595_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_596_root_address_inst
    process(array_obj_ref_596_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_596_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_596_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_811_index_2_rename
    process(R_ix_x1293_810_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1293_810_resized;
      ov(14 downto 0) := iv;
      R_ix_x1293_810_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_811_index_2_resize
    process(ix_x1293_797) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1293_797;
      ov := iv(14 downto 0);
      R_ix_x1293_810_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_811_root_address_inst
    process(array_obj_ref_811_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_811_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_811_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1041_addr_0
    process(ptr_deref_1041_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1041_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_1041_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1041_base_resize
    process(arrayidx219_1038) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx219_1038;
      ov := iv(14 downto 0);
      ptr_deref_1041_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1041_gather_scatter
    process(ptr_deref_1041_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1041_data_0;
      ov(63 downto 0) := iv;
      tmp220_1042 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1041_root_address_inst
    process(ptr_deref_1041_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1041_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_1041_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_733_addr_0
    process(ptr_deref_733_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_733_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_733_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_733_base_resize
    process(arrayidx_598) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_598;
      ov := iv(14 downto 0);
      ptr_deref_733_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_733_gather_scatter
    process(add115_731) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add115_731;
      ov(63 downto 0) := iv;
      ptr_deref_733_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_733_root_address_inst
    process(ptr_deref_733_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_733_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_733_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_815_addr_0
    process(ptr_deref_815_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_815_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_815_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_815_base_resize
    process(arrayidx127_813) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx127_813;
      ov := iv(14 downto 0);
      ptr_deref_815_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_815_gather_scatter
    process(type_cast_817_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_817_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_815_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_815_root_address_inst
    process(ptr_deref_815_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_815_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_815_root_address <= ov(14 downto 0);
      --
    end process;
    if_stmt_1152_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond8_1151;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1152_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1152_branch_req_0,
          ack0 => if_stmt_1152_branch_ack_0,
          ack1 => if_stmt_1152_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_517_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp296_516;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_517_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_517_branch_req_0,
          ack0 => if_stmt_517_branch_ack_0,
          ack1 => if_stmt_517_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_532_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp123292_531;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_532_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_532_branch_req_0,
          ack0 => if_stmt_532_branch_ack_0,
          ack1 => if_stmt_532_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_747_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond24_746;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_747_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_747_branch_req_0,
          ack0 => if_stmt_747_branch_ack_0,
          ack1 => if_stmt_747_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_830_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_829;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_830_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_830_branch_req_0,
          ack0 => if_stmt_830_branch_ack_0,
          ack1 => if_stmt_830_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_972_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp123292_531;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_972_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_972_branch_req_0,
          ack0 => if_stmt_972_branch_ack_0,
          ack1 => if_stmt_972_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1145_inst
    process(ix_x2290_1022) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x2290_1022, type_cast_1144_wire_constant, tmp_var);
      inc286_1146 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_740_inst
    process(ix_x0297_582) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x0297_582, type_cast_739_wire_constant, tmp_var);
      inc_741 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_823_inst
    process(ix_x1293_797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x1293_797, type_cast_822_wire_constant, tmp_var);
      inc130_824 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1150_inst
    process(inc286_1146, umax7_1019) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc286_1146, umax7_1019, tmp_var);
      exitcond8_1151 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_745_inst
    process(inc_741, umax23_579) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_741, umax23_579, tmp_var);
      exitcond24_746 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_828_inst
    process(inc130_824, umax_794) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc130_824, umax_794, tmp_var);
      exitcond_829 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1005_inst
    process(tmp4_1000) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1000, type_cast_1004_wire_constant, tmp_var);
      tmp5_1006 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_565_inst
    process(tmp20_560) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_560, type_cast_564_wire_constant, tmp_var);
      tmp21_566 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_780_inst
    process(tmp13_775) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp13_775, type_cast_779_wire_constant, tmp_var);
      tmp14_781 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1051_inst
    process(tmp220_1042) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp220_1042, type_cast_1050_wire_constant, tmp_var);
      shr227_1052 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1061_inst
    process(tmp220_1042) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp220_1042, type_cast_1060_wire_constant, tmp_var);
      shr233_1062 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1071_inst
    process(tmp220_1042) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp220_1042, type_cast_1070_wire_constant, tmp_var);
      shr239_1072 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1081_inst
    process(tmp220_1042) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp220_1042, type_cast_1080_wire_constant, tmp_var);
      shr245_1082 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1091_inst
    process(tmp220_1042) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp220_1042, type_cast_1090_wire_constant, tmp_var);
      shr251_1092 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1101_inst
    process(tmp220_1042) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp220_1042, type_cast_1100_wire_constant, tmp_var);
      shr257_1102 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1111_inst
    process(tmp220_1042) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp220_1042, type_cast_1110_wire_constant, tmp_var);
      shr263_1112 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_881_inst
    process(sub_872) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_872, type_cast_880_wire_constant, tmp_var);
      shr152_882 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_891_inst
    process(sub_872) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_872, type_cast_890_wire_constant, tmp_var);
      shr158_892 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_901_inst
    process(sub_872) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_872, type_cast_900_wire_constant, tmp_var);
      shr164_902 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_911_inst
    process(sub_872) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_872, type_cast_910_wire_constant, tmp_var);
      shr170_912 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_921_inst
    process(sub_872) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_872, type_cast_920_wire_constant, tmp_var);
      shr176_922 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_931_inst
    process(sub_872) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_872, type_cast_930_wire_constant, tmp_var);
      shr182_932 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_941_inst
    process(sub_872) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_872, type_cast_940_wire_constant, tmp_var);
      shr188_942 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_482_inst
    process(conv55_474, conv53_470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv55_474, conv53_470, tmp_var);
      mul_483 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_487_inst
    process(mul_483, conv57_478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_483, conv57_478, tmp_var);
      mul58_488 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_504_inst
    process(conv63_496, conv61_492) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_496, conv61_492, tmp_var);
      mul64_505 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_509_inst
    process(mul64_505, conv66_500) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul64_505, conv66_500, tmp_var);
      mul67_510 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_550_inst
    process(tmp16_542, tmp17_546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_542, tmp17_546, tmp_var);
      tmp18_551 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_559_inst
    process(tmp18_551, tmp19_555) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp18_551, tmp19_555, tmp_var);
      tmp20_560 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_765_inst
    process(tmp9_757, tmp10_761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_757, tmp10_761, tmp_var);
      tmp11_766 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_774_inst
    process(tmp11_766, tmp12_770) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp11_766, tmp12_770, tmp_var);
      tmp13_775 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_990_inst
    process(tmp_982, tmp1_986) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_982, tmp1_986, tmp_var);
      tmp2_991 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_999_inst
    process(tmp2_991, tmp3_995) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_991, tmp3_995, tmp_var);
      tmp4_1000 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_340_inst
    process(shl_329, conv3_336) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_329, conv3_336, tmp_var);
      add_341 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_365_inst
    process(shl9_354, conv11_361) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_354, conv11_361, tmp_var);
      add12_366 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_390_inst
    process(shl18_379, conv20_386) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_379, conv20_386, tmp_var);
      add21_391 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_415_inst
    process(shl27_404, conv29_411) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_404, conv29_411, tmp_var);
      add30_416 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_440_inst
    process(shl36_429, conv38_436) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_429, conv38_436, tmp_var);
      add39_441 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_465_inst
    process(shl45_454, conv47_461) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_454, conv47_461, tmp_var);
      add48_466 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_622_inst
    process(shl75_611, conv78_618) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl75_611, conv78_618, tmp_var);
      add79_623 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_640_inst
    process(shl81_629, conv84_636) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl81_629, conv84_636, tmp_var);
      add85_641 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_658_inst
    process(shl87_647, conv90_654) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl87_647, conv90_654, tmp_var);
      add91_659 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_676_inst
    process(shl93_665, conv96_672) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl93_665, conv96_672, tmp_var);
      add97_677 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_694_inst
    process(shl99_683, conv102_690) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl99_683, conv102_690, tmp_var);
      add103_695 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_712_inst
    process(shl105_701, conv108_708) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_701, conv108_708, tmp_var);
      add109_713 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_730_inst
    process(shl111_719, conv114_726) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl111_719, conv114_726, tmp_var);
      add115_731 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_328_inst
    process(conv1_323) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_323, type_cast_327_wire_constant, tmp_var);
      shl_329 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_353_inst
    process(conv8_348) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_348, type_cast_352_wire_constant, tmp_var);
      shl9_354 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_378_inst
    process(conv17_373) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_373, type_cast_377_wire_constant, tmp_var);
      shl18_379 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_403_inst
    process(conv26_398) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_398, type_cast_402_wire_constant, tmp_var);
      shl27_404 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_428_inst
    process(conv35_423) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_423, type_cast_427_wire_constant, tmp_var);
      shl36_429 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_453_inst
    process(conv44_448) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_448, type_cast_452_wire_constant, tmp_var);
      shl45_454 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_610_inst
    process(conv73_605) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv73_605, type_cast_609_wire_constant, tmp_var);
      shl75_611 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_628_inst
    process(add79_623) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add79_623, type_cast_627_wire_constant, tmp_var);
      shl81_629 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_646_inst
    process(add85_641) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add85_641, type_cast_645_wire_constant, tmp_var);
      shl87_647 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_664_inst
    process(add91_659) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add91_659, type_cast_663_wire_constant, tmp_var);
      shl93_665 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_682_inst
    process(add97_677) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add97_677, type_cast_681_wire_constant, tmp_var);
      shl99_683 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_700_inst
    process(add103_695) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add103_695, type_cast_699_wire_constant, tmp_var);
      shl105_701 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_718_inst
    process(add109_713) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add109_713, type_cast_717_wire_constant, tmp_var);
      shl111_719 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_871_inst
    process(conv143_867, conv134_847) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv143_867, conv134_847, tmp_var);
      sub_872 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1011_inst
    process(tmp5_1006) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp5_1006, type_cast_1010_wire_constant, tmp_var);
      tmp6_1012 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_515_inst
    process(mul58_488) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul58_488, type_cast_514_wire_constant, tmp_var);
      cmp296_516 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_530_inst
    process(mul67_510) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul67_510, type_cast_529_wire_constant, tmp_var);
      cmp123292_531 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_571_inst
    process(tmp21_566) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp21_566, type_cast_570_wire_constant, tmp_var);
      tmp22_572 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_786_inst
    process(tmp14_781) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp14_781, type_cast_785_wire_constant, tmp_var);
      tmp15_787 <= tmp_var; --
    end process;
    -- shared split operator group (65) : array_obj_ref_1036_index_offset 
    ApIntAdd_group_65: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x2290_1035_scaled;
      array_obj_ref_1036_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1036_index_offset_req_0;
      array_obj_ref_1036_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1036_index_offset_req_1;
      array_obj_ref_1036_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_65_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_65_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "100000000000000",
          constant_width => 15,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : array_obj_ref_596_index_offset 
    ApIntAdd_group_66: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0297_595_scaled;
      array_obj_ref_596_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_596_index_offset_req_0;
      array_obj_ref_596_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_596_index_offset_req_1;
      array_obj_ref_596_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_66_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_66_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "000000000000000",
          constant_width => 15,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : array_obj_ref_811_index_offset 
    ApIntAdd_group_67: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1293_810_scaled;
      array_obj_ref_811_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_811_index_offset_req_0;
      array_obj_ref_811_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_811_index_offset_req_1;
      array_obj_ref_811_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_67_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_67_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_67",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "100000000000000",
          constant_width => 15,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- unary operator type_cast_845_inst
    process(call133_841) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call133_841, tmp_var);
      type_cast_845_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_865_inst
    process(call142_862) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call142_862, tmp_var);
      type_cast_865_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1041_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1041_load_0_req_0;
      ptr_deref_1041_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1041_load_0_req_1;
      ptr_deref_1041_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1041_word_address_0;
      ptr_deref_1041_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 15,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(14 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_815_store_0 ptr_deref_733_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(29 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_815_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_733_store_0_req_0;
      ptr_deref_815_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_733_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_815_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_733_store_0_req_1;
      ptr_deref_815_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_733_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_815_word_address_0 & ptr_deref_733_word_address_0;
      data_in <= ptr_deref_815_data_0 & ptr_deref_733_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 15,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(14 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Zeropad_input_pipe_318_inst RPIPE_Zeropad_input_pipe_331_inst RPIPE_Zeropad_input_pipe_343_inst RPIPE_Zeropad_input_pipe_356_inst RPIPE_Zeropad_input_pipe_368_inst RPIPE_Zeropad_input_pipe_381_inst RPIPE_Zeropad_input_pipe_393_inst RPIPE_Zeropad_input_pipe_406_inst RPIPE_Zeropad_input_pipe_418_inst RPIPE_Zeropad_input_pipe_431_inst RPIPE_Zeropad_input_pipe_443_inst RPIPE_Zeropad_input_pipe_456_inst RPIPE_Zeropad_input_pipe_600_inst RPIPE_Zeropad_input_pipe_613_inst RPIPE_Zeropad_input_pipe_631_inst RPIPE_Zeropad_input_pipe_649_inst RPIPE_Zeropad_input_pipe_667_inst RPIPE_Zeropad_input_pipe_685_inst RPIPE_Zeropad_input_pipe_703_inst RPIPE_Zeropad_input_pipe_721_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(159 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 19 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 19 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 19 downto 0);
      signal guard_vector : std_logic_vector( 19 downto 0);
      constant outBUFs : IntegerArray(19 downto 0) := (19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(19 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false);
      constant guardBuffering: IntegerArray(19 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2);
      -- 
    begin -- 
      reqL_unguarded(19) <= RPIPE_Zeropad_input_pipe_318_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Zeropad_input_pipe_331_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Zeropad_input_pipe_343_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Zeropad_input_pipe_356_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Zeropad_input_pipe_368_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Zeropad_input_pipe_381_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Zeropad_input_pipe_393_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Zeropad_input_pipe_406_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Zeropad_input_pipe_418_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Zeropad_input_pipe_431_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Zeropad_input_pipe_443_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Zeropad_input_pipe_456_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Zeropad_input_pipe_600_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Zeropad_input_pipe_613_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Zeropad_input_pipe_631_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Zeropad_input_pipe_649_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Zeropad_input_pipe_667_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Zeropad_input_pipe_685_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Zeropad_input_pipe_703_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Zeropad_input_pipe_721_inst_req_0;
      RPIPE_Zeropad_input_pipe_318_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Zeropad_input_pipe_331_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Zeropad_input_pipe_343_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Zeropad_input_pipe_356_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Zeropad_input_pipe_368_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Zeropad_input_pipe_381_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Zeropad_input_pipe_393_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Zeropad_input_pipe_406_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Zeropad_input_pipe_418_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Zeropad_input_pipe_431_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Zeropad_input_pipe_443_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Zeropad_input_pipe_456_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Zeropad_input_pipe_600_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Zeropad_input_pipe_613_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Zeropad_input_pipe_631_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Zeropad_input_pipe_649_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Zeropad_input_pipe_667_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Zeropad_input_pipe_685_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Zeropad_input_pipe_703_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Zeropad_input_pipe_721_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(19) <= RPIPE_Zeropad_input_pipe_318_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Zeropad_input_pipe_331_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Zeropad_input_pipe_343_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Zeropad_input_pipe_356_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Zeropad_input_pipe_368_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Zeropad_input_pipe_381_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Zeropad_input_pipe_393_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Zeropad_input_pipe_406_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Zeropad_input_pipe_418_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Zeropad_input_pipe_431_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Zeropad_input_pipe_443_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Zeropad_input_pipe_456_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Zeropad_input_pipe_600_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Zeropad_input_pipe_613_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Zeropad_input_pipe_631_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Zeropad_input_pipe_649_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Zeropad_input_pipe_667_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Zeropad_input_pipe_685_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Zeropad_input_pipe_703_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Zeropad_input_pipe_721_inst_req_1;
      RPIPE_Zeropad_input_pipe_318_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Zeropad_input_pipe_331_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Zeropad_input_pipe_343_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Zeropad_input_pipe_356_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Zeropad_input_pipe_368_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Zeropad_input_pipe_381_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Zeropad_input_pipe_393_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Zeropad_input_pipe_406_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Zeropad_input_pipe_418_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Zeropad_input_pipe_431_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Zeropad_input_pipe_443_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Zeropad_input_pipe_456_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Zeropad_input_pipe_600_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Zeropad_input_pipe_613_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Zeropad_input_pipe_631_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Zeropad_input_pipe_649_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Zeropad_input_pipe_667_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Zeropad_input_pipe_685_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Zeropad_input_pipe_703_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Zeropad_input_pipe_721_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      call_319 <= data_out(159 downto 152);
      call2_332 <= data_out(151 downto 144);
      call5_344 <= data_out(143 downto 136);
      call10_357 <= data_out(135 downto 128);
      call14_369 <= data_out(127 downto 120);
      call19_382 <= data_out(119 downto 112);
      call23_394 <= data_out(111 downto 104);
      call28_407 <= data_out(103 downto 96);
      call32_419 <= data_out(95 downto 88);
      call37_432 <= data_out(87 downto 80);
      call41_444 <= data_out(79 downto 72);
      call46_457 <= data_out(71 downto 64);
      call72_601 <= data_out(63 downto 56);
      call76_614 <= data_out(55 downto 48);
      call82_632 <= data_out(47 downto 40);
      call88_650 <= data_out(39 downto 32);
      call94_668 <= data_out(31 downto 24);
      call100_686 <= data_out(23 downto 16);
      call106_704 <= data_out(15 downto 8);
      call112_722 <= data_out(7 downto 0);
      Zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "Zeropad_input_pipe_read_0_gI", nreqs => 20, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "Zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 20,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Zeropad_input_pipe_pipe_read_req(0),
          oack => Zeropad_input_pipe_pipe_read_ack(0),
          odata => Zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Zeropad_output_pipe_1123_inst WPIPE_Zeropad_output_pipe_1135_inst WPIPE_Zeropad_output_pipe_1138_inst WPIPE_Zeropad_output_pipe_1126_inst WPIPE_Zeropad_output_pipe_1129_inst WPIPE_Zeropad_output_pipe_947_inst WPIPE_Zeropad_output_pipe_950_inst WPIPE_Zeropad_output_pipe_1120_inst WPIPE_Zeropad_output_pipe_1132_inst WPIPE_Zeropad_output_pipe_953_inst WPIPE_Zeropad_output_pipe_956_inst WPIPE_Zeropad_output_pipe_1117_inst WPIPE_Zeropad_output_pipe_959_inst WPIPE_Zeropad_output_pipe_962_inst WPIPE_Zeropad_output_pipe_965_inst WPIPE_Zeropad_output_pipe_968_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_Zeropad_output_pipe_1123_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Zeropad_output_pipe_1135_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Zeropad_output_pipe_1138_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Zeropad_output_pipe_1126_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Zeropad_output_pipe_1129_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Zeropad_output_pipe_947_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Zeropad_output_pipe_950_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Zeropad_output_pipe_1120_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Zeropad_output_pipe_1132_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Zeropad_output_pipe_953_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Zeropad_output_pipe_956_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Zeropad_output_pipe_1117_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Zeropad_output_pipe_959_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Zeropad_output_pipe_962_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Zeropad_output_pipe_965_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Zeropad_output_pipe_968_inst_req_0;
      WPIPE_Zeropad_output_pipe_1123_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Zeropad_output_pipe_1135_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Zeropad_output_pipe_1138_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Zeropad_output_pipe_1126_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Zeropad_output_pipe_1129_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Zeropad_output_pipe_947_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Zeropad_output_pipe_950_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Zeropad_output_pipe_1120_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Zeropad_output_pipe_1132_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Zeropad_output_pipe_953_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Zeropad_output_pipe_956_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Zeropad_output_pipe_1117_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Zeropad_output_pipe_959_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Zeropad_output_pipe_962_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Zeropad_output_pipe_965_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Zeropad_output_pipe_968_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_Zeropad_output_pipe_1123_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Zeropad_output_pipe_1135_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Zeropad_output_pipe_1138_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Zeropad_output_pipe_1126_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Zeropad_output_pipe_1129_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Zeropad_output_pipe_947_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Zeropad_output_pipe_950_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Zeropad_output_pipe_1120_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Zeropad_output_pipe_1132_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Zeropad_output_pipe_953_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Zeropad_output_pipe_956_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Zeropad_output_pipe_1117_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Zeropad_output_pipe_959_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Zeropad_output_pipe_962_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Zeropad_output_pipe_965_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Zeropad_output_pipe_968_inst_req_1;
      WPIPE_Zeropad_output_pipe_1123_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Zeropad_output_pipe_1135_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Zeropad_output_pipe_1138_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Zeropad_output_pipe_1126_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Zeropad_output_pipe_1129_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Zeropad_output_pipe_947_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Zeropad_output_pipe_950_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Zeropad_output_pipe_1120_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Zeropad_output_pipe_1132_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Zeropad_output_pipe_953_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Zeropad_output_pipe_956_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Zeropad_output_pipe_1117_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Zeropad_output_pipe_959_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Zeropad_output_pipe_962_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Zeropad_output_pipe_965_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Zeropad_output_pipe_968_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv254_1096 & conv230_1056 & conv224_1046 & conv248_1086 & conv242_1076 & conv191_946 & conv185_936 & conv260_1106 & conv236_1066 & conv179_926 & conv173_916 & conv266_1116 & conv167_906 & conv161_896 & conv155_886 & conv149_876;
      Zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "Zeropad_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "Zeropad_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Zeropad_output_pipe_pipe_write_req(0),
          oack => Zeropad_output_pipe_pipe_write_ack(0),
          odata => Zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_841_call call_stmt_862_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_841_call_req_0;
      reqL_unguarded(0) <= call_stmt_862_call_req_0;
      call_stmt_841_call_ack_0 <= ackL_unguarded(1);
      call_stmt_862_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_841_call_req_1;
      reqR_unguarded(0) <= call_stmt_862_call_req_1;
      call_stmt_841_call_ack_1 <= ackR_unguarded(1);
      call_stmt_862_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call133_841 <= data_out(127 downto 64);
      call142_862 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_859_call 
    zeropad_same_call_group_1: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_859_call_req_0;
      call_stmt_859_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_859_call_req_1;
      call_stmt_859_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      zeropad_same_call_group_1_gI: SplitGuardInterface generic map(name => "zeropad_same_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add_341 & add12_366 & add21_391 & add30_416 & add39_441 & add48_466 & type_cast_856_wire_constant & type_cast_858_wire_constant;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 112,
        owidth => 112,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => zeropad_same_call_reqs(0),
          ackR => zeropad_same_call_acks(0),
          dataR => zeropad_same_call_data(111 downto 0),
          tagR => zeropad_same_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => zeropad_same_return_acks(0), -- cross-over
          ackL => zeropad_same_return_reqs(0), -- cross-over
          tagL => zeropad_same_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad_same is -- 
  generic (tag_length : integer); 
  port ( -- 
    inp_d0 : in  std_logic_vector(15 downto 0);
    inp_d1 : in  std_logic_vector(15 downto 0);
    inp_d2 : in  std_logic_vector(15 downto 0);
    out_d0 : in  std_logic_vector(15 downto 0);
    out_d1 : in  std_logic_vector(15 downto 0);
    out_d2 : in  std_logic_vector(15 downto 0);
    index1 : in  std_logic_vector(7 downto 0);
    index2 : in  std_logic_vector(7 downto 0);
    readModule1_call_reqs : out  std_logic_vector(0 downto 0);
    readModule1_call_acks : in   std_logic_vector(0 downto 0);
    readModule1_call_data : out  std_logic_vector(39 downto 0);
    readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
    readModule1_return_reqs : out  std_logic_vector(0 downto 0);
    readModule1_return_acks : in   std_logic_vector(0 downto 0);
    readModule1_return_data : in   std_logic_vector(63 downto 0);
    readModule1_return_tag :  in   std_logic_vector(0 downto 0);
    writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
    writeModule1_call_acks : in   std_logic_vector(0 downto 0);
    writeModule1_call_data : out  std_logic_vector(103 downto 0);
    writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
    writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
    writeModule1_return_acks : in   std_logic_vector(0 downto 0);
    writeModule1_return_data : in   std_logic_vector(0 downto 0);
    writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad_same;
architecture zeropad_same_arch of zeropad_same is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 112)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal inp_d0_buffer :  std_logic_vector(15 downto 0);
  signal inp_d0_update_enable: Boolean;
  signal inp_d1_buffer :  std_logic_vector(15 downto 0);
  signal inp_d1_update_enable: Boolean;
  signal inp_d2_buffer :  std_logic_vector(15 downto 0);
  signal inp_d2_update_enable: Boolean;
  signal out_d0_buffer :  std_logic_vector(15 downto 0);
  signal out_d0_update_enable: Boolean;
  signal out_d1_buffer :  std_logic_vector(15 downto 0);
  signal out_d1_update_enable: Boolean;
  signal out_d2_buffer :  std_logic_vector(15 downto 0);
  signal out_d2_update_enable: Boolean;
  signal index1_buffer :  std_logic_vector(7 downto 0);
  signal index1_update_enable: Boolean;
  signal index2_buffer :  std_logic_vector(7 downto 0);
  signal index2_update_enable: Boolean;
  -- output port buffer signals
  signal zeropad_same_CP_493_start: Boolean;
  signal zeropad_same_CP_493_symbol: Boolean;
  -- volatile/operator module components. 
  component readModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(14 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      done : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(14 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal phi_stmt_132_ack_0 : boolean;
  signal next_add_dest_dim0_272_143_buf_ack_0 : boolean;
  signal add_dest_dim0_init_118_142_buf_ack_0 : boolean;
  signal add_dest_dim0_init_118_142_buf_ack_1 : boolean;
  signal phi_stmt_128_req_0 : boolean;
  signal add_dest_dim0_init_118_142_buf_req_1 : boolean;
  signal next_add_dest_dim1_266_146_buf_ack_1 : boolean;
  signal next_add_dest_dim1_266_146_buf_ack_0 : boolean;
  signal phi_stmt_128_req_1 : boolean;
  signal next_input_dim2_278_139_buf_req_0 : boolean;
  signal add_dest_dim1_init_121_147_buf_req_0 : boolean;
  signal add_dest_dim0_init_118_142_buf_req_0 : boolean;
  signal phi_stmt_140_req_0 : boolean;
  signal add_dest_dim1_init_121_147_buf_ack_0 : boolean;
  signal phi_stmt_140_req_1 : boolean;
  signal next_add_dest_dim1_266_146_buf_req_0 : boolean;
  signal next_add_dest_dim0_272_143_buf_req_0 : boolean;
  signal phi_stmt_148_req_1 : boolean;
  signal next_add_dest_dim0_272_143_buf_ack_1 : boolean;
  signal next_add_dest_dim1_266_146_buf_req_1 : boolean;
  signal call_stmt_182_call_req_0 : boolean;
  signal call_stmt_182_call_ack_0 : boolean;
  signal type_cast_185_inst_req_0 : boolean;
  signal type_cast_185_inst_ack_0 : boolean;
  signal next_add_src_253_151_buf_ack_0 : boolean;
  signal call_stmt_191_call_req_1 : boolean;
  signal call_stmt_191_call_ack_1 : boolean;
  signal next_input_dim0_294_131_buf_ack_0 : boolean;
  signal phi_stmt_144_req_0 : boolean;
  signal next_input_dim0_294_131_buf_req_0 : boolean;
  signal next_input_dim2_278_139_buf_ack_1 : boolean;
  signal phi_stmt_136_req_0 : boolean;
  signal phi_stmt_132_req_0 : boolean;
  signal next_input_dim1_288_135_buf_ack_1 : boolean;
  signal next_input_dim1_288_135_buf_req_1 : boolean;
  signal add_dest_dim1_init_121_147_buf_ack_1 : boolean;
  signal next_input_dim1_288_135_buf_ack_0 : boolean;
  signal next_add_dest_dim0_272_143_buf_req_1 : boolean;
  signal next_input_dim2_278_139_buf_req_1 : boolean;
  signal next_input_dim1_288_135_buf_req_0 : boolean;
  signal phi_stmt_132_req_1 : boolean;
  signal phi_stmt_140_ack_0 : boolean;
  signal next_add_src_253_151_buf_req_1 : boolean;
  signal call_stmt_182_call_req_1 : boolean;
  signal call_stmt_182_call_ack_1 : boolean;
  signal phi_stmt_136_ack_0 : boolean;
  signal call_stmt_191_call_req_0 : boolean;
  signal call_stmt_191_call_ack_0 : boolean;
  signal do_while_stmt_126_branch_req_0 : boolean;
  signal next_input_dim2_278_139_buf_ack_0 : boolean;
  signal next_input_dim0_294_131_buf_ack_1 : boolean;
  signal next_input_dim0_294_131_buf_req_1 : boolean;
  signal phi_stmt_128_ack_0 : boolean;
  signal phi_stmt_136_req_1 : boolean;
  signal next_add_src_253_151_buf_req_0 : boolean;
  signal phi_stmt_148_ack_0 : boolean;
  signal phi_stmt_148_req_0 : boolean;
  signal add_dest_dim1_init_121_147_buf_req_1 : boolean;
  signal phi_stmt_144_req_1 : boolean;
  signal next_add_src_253_151_buf_ack_1 : boolean;
  signal type_cast_185_inst_req_1 : boolean;
  signal type_cast_185_inst_ack_1 : boolean;
  signal phi_stmt_144_ack_0 : boolean;
  signal W_dim2_limit_196_delayed_1_0_197_inst_req_0 : boolean;
  signal W_dim2_limit_196_delayed_1_0_197_inst_ack_0 : boolean;
  signal W_dim2_limit_196_delayed_1_0_197_inst_req_1 : boolean;
  signal W_dim2_limit_196_delayed_1_0_197_inst_ack_1 : boolean;
  signal SUB_u16_u16_208_inst_req_0 : boolean;
  signal SUB_u16_u16_208_inst_ack_0 : boolean;
  signal SUB_u16_u16_208_inst_req_1 : boolean;
  signal SUB_u16_u16_208_inst_ack_1 : boolean;
  signal W_nid1_true4_249_delayed_1_0_254_inst_req_0 : boolean;
  signal W_nid1_true4_249_delayed_1_0_254_inst_ack_0 : boolean;
  signal W_nid1_true4_249_delayed_1_0_254_inst_req_1 : boolean;
  signal W_nid1_true4_249_delayed_1_0_254_inst_ack_1 : boolean;
  signal SUB_u16_u16_298_inst_req_0 : boolean;
  signal SUB_u16_u16_298_inst_ack_0 : boolean;
  signal SUB_u16_u16_298_inst_req_1 : boolean;
  signal SUB_u16_u16_298_inst_ack_1 : boolean;
  signal do_while_stmt_126_branch_ack_0 : boolean;
  signal do_while_stmt_126_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad_same_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 112) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= inp_d0;
  inp_d0_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= inp_d1;
  inp_d1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= inp_d2;
  inp_d2_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= out_d0;
  out_d0_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= out_d1;
  out_d1_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= out_d2;
  out_d2_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(103 downto 96) <= index1;
  index1_buffer <= in_buffer_data_out(103 downto 96);
  in_buffer_data_in(111 downto 104) <= index2;
  index2_buffer <= in_buffer_data_out(111 downto 104);
  in_buffer_data_in(tag_length + 111 downto 112) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 111 downto 112);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad_same_CP_493_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad_same_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad_same_CP_493_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad_same_CP_493_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad_same_CP_493_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad_same_CP_493: Block -- control-path 
    signal zeropad_same_CP_493_elements: BooleanArray(159 downto 0);
    -- 
  begin -- 
    zeropad_same_CP_493_elements(0) <= zeropad_same_CP_493_start;
    zeropad_same_CP_493_symbol <= zeropad_same_CP_493_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_96/do_while_stmt_126__entry__
      -- CP-element group 0: 	 branch_block_stmt_96/assign_stmt_100_to_assign_stmt_125__exit__
      -- CP-element group 0: 	 branch_block_stmt_96/assign_stmt_100_to_assign_stmt_125__entry__
      -- CP-element group 0: 	 branch_block_stmt_96/assign_stmt_100_to_assign_stmt_125/$exit
      -- CP-element group 0: 	 branch_block_stmt_96/assign_stmt_100_to_assign_stmt_125/$entry
      -- CP-element group 0: 	 branch_block_stmt_96/branch_block_stmt_96__entry__
      -- CP-element group 0: 	 branch_block_stmt_96/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	159 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_96/do_while_stmt_126__exit__
      -- CP-element group 1: 	 branch_block_stmt_96/branch_block_stmt_96__exit__
      -- CP-element group 1: 	 branch_block_stmt_96/$exit
      -- 
    zeropad_same_CP_493_elements(1) <= zeropad_same_CP_493_elements(159);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126__entry__
      -- CP-element group 2: 	 branch_block_stmt_96/do_while_stmt_126/$entry
      -- 
    zeropad_same_CP_493_elements(2) <= zeropad_same_CP_493_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	159 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126__exit__
      -- 
    -- Element group zeropad_same_CP_493_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_96/do_while_stmt_126/loop_back
      -- 
    -- Element group zeropad_same_CP_493_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	157 
    -- CP-element group 5: 	158 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_96/do_while_stmt_126/condition_done
      -- CP-element group 5: 	 branch_block_stmt_96/do_while_stmt_126/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_96/do_while_stmt_126/loop_taken/$entry
      -- 
    zeropad_same_CP_493_elements(5) <= zeropad_same_CP_493_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	156 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_96/do_while_stmt_126/loop_body_done
      -- 
    zeropad_same_CP_493_elements(6) <= zeropad_same_CP_493_elements(156);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	95 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	114 
    -- CP-element group 7: 	59 
    -- CP-element group 7: 	78 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/back_edge_to_loop_body
      -- 
    zeropad_same_CP_493_elements(7) <= zeropad_same_CP_493_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	97 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	116 
    -- CP-element group 8: 	61 
    -- CP-element group 8: 	80 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/first_time_through_loop_body
      -- 
    zeropad_same_CP_493_elements(8) <= zeropad_same_CP_493_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	91 
    -- CP-element group 9: 	92 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	108 
    -- CP-element group 9: 	109 
    -- CP-element group 9: 	139 
    -- CP-element group 9: 	143 
    -- CP-element group 9: 	155 
    -- CP-element group 9: 	147 
    -- CP-element group 9: 	151 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	54 
    -- CP-element group 9: 	72 
    -- CP-element group 9: 	73 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/loop_body_start
      -- 
    -- Element group zeropad_same_CP_493_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	142 
    -- CP-element group 10: 	154 
    -- CP-element group 10: 	155 
    -- CP-element group 10: 	146 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/condition_evaluated
      -- 
    condition_evaluated_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(10), ack => do_while_stmt_126_branch_req_0); -- 
    zeropad_same_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(14) & zeropad_same_CP_493_elements(142) & zeropad_same_CP_493_elements(154) & zeropad_same_CP_493_elements(155) & zeropad_same_CP_493_elements(146);
      gj_zeropad_same_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	91 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	108 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	110 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	74 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/aggregated_phi_sample_req
      -- 
    zeropad_same_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(91) & zeropad_same_CP_493_elements(15) & zeropad_same_CP_493_elements(34) & zeropad_same_CP_493_elements(108) & zeropad_same_CP_493_elements(53) & zeropad_same_CP_493_elements(72) & zeropad_same_CP_493_elements(14);
      gj_zeropad_same_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	93 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	111 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	75 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	140 
    -- CP-element group 12: 	144 
    -- CP-element group 12: 	156 
    -- CP-element group 12: 	148 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	91 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	108 
    -- CP-element group 12: 	53 
    -- CP-element group 12: 	72 
    -- CP-element group 12:  members (7) 
      -- CP-element group 12: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_sample_completed_
      -- 
    zeropad_same_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(93) & zeropad_same_CP_493_elements(18) & zeropad_same_CP_493_elements(37) & zeropad_same_CP_493_elements(111) & zeropad_same_CP_493_elements(56) & zeropad_same_CP_493_elements(75);
      gj_zeropad_same_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	92 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	109 
    -- CP-element group 13: 	54 
    -- CP-element group 13: 	73 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	112 
    -- CP-element group 13: 	57 
    -- CP-element group 13: 	76 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/aggregated_phi_update_req
      -- 
    zeropad_same_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(92) & zeropad_same_CP_493_elements(16) & zeropad_same_CP_493_elements(35) & zeropad_same_CP_493_elements(109) & zeropad_same_CP_493_elements(54) & zeropad_same_CP_493_elements(73);
      gj_zeropad_same_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	94 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	113 
    -- CP-element group 14: 	58 
    -- CP-element group 14: 	77 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/aggregated_phi_update_ack
      -- 
    zeropad_same_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(94) & zeropad_same_CP_493_elements(20) & zeropad_same_CP_493_elements(39) & zeropad_same_CP_493_elements(113) & zeropad_same_CP_493_elements(58) & zeropad_same_CP_493_elements(77);
      gj_zeropad_same_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: 	142 
    -- CP-element group 15: 	146 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_sample_start_
      -- 
    zeropad_same_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(142) & zeropad_same_CP_493_elements(146);
      gj_zeropad_same_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_update_start_
      -- 
    zeropad_same_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(20);
      gj_zeropad_same_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_sample_start__ps
      -- 
    zeropad_same_CP_493_elements(17) <= zeropad_same_CP_493_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_update_start__ps
      -- 
    zeropad_same_CP_493_elements(19) <= zeropad_same_CP_493_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_loopback_trigger
      -- 
    zeropad_same_CP_493_elements(21) <= zeropad_same_CP_493_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_loopback_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_loopback_sample_req
      -- 
    phi_stmt_128_loopback_sample_req_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_128_loopback_sample_req_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(22), ack => phi_stmt_128_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_entry_trigger
      -- 
    zeropad_same_CP_493_elements(23) <= zeropad_same_CP_493_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_entry_sample_req_ps
      -- CP-element group 24: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_entry_sample_req
      -- 
    phi_stmt_128_entry_sample_req_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_128_entry_sample_req_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(24), ack => phi_stmt_128_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_phi_mux_ack_ps
      -- CP-element group 25: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_128_phi_mux_ack
      -- 
    phi_stmt_128_phi_mux_ack_543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_128_ack_0, ack => zeropad_same_CP_493_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim0_init_130_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim0_init_130_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim0_init_130_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim0_init_130_sample_start_
      -- 
    -- Element group zeropad_same_CP_493_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim0_init_130_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim0_init_130_update_start_
      -- 
    -- Element group zeropad_same_CP_493_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim0_init_130_update_completed__ps
      -- 
    zeropad_same_CP_493_elements(28) <= zeropad_same_CP_493_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim0_init_130_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => zeropad_same_CP_493_elements(27), ack => zeropad_same_CP_493_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_Sample/req
      -- CP-element group 30: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_Sample/$entry
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(30), ack => next_input_dim0_294_131_buf_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_update_start_
      -- CP-element group 31: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_Update/req
      -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(31), ack => next_input_dim0_294_131_buf_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_Sample/ack
      -- CP-element group 32: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_sample_completed_
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim0_294_131_buf_ack_0, ack => zeropad_same_CP_493_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim0_131_Update/ack
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim0_294_131_buf_ack_1, ack => zeropad_same_CP_493_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: 	142 
    -- CP-element group 34: 	146 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_sample_start_
      -- 
    zeropad_same_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(142) & zeropad_same_CP_493_elements(146);
      gj_zeropad_same_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	39 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_update_start_
      -- 
    zeropad_same_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(39);
      gj_zeropad_same_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_sample_start__ps
      -- 
    zeropad_same_CP_493_elements(36) <= zeropad_same_CP_493_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_update_start__ps
      -- 
    zeropad_same_CP_493_elements(38) <= zeropad_same_CP_493_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	35 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_update_completed__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_loopback_trigger
      -- 
    zeropad_same_CP_493_elements(40) <= zeropad_same_CP_493_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_loopback_sample_req_ps
      -- CP-element group 41: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_loopback_sample_req
      -- 
    phi_stmt_132_loopback_sample_req_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_132_loopback_sample_req_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(41), ack => phi_stmt_132_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_entry_trigger
      -- 
    zeropad_same_CP_493_elements(42) <= zeropad_same_CP_493_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_entry_sample_req_ps
      -- CP-element group 43: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_entry_sample_req
      -- 
    phi_stmt_132_entry_sample_req_584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_132_entry_sample_req_584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(43), ack => phi_stmt_132_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_132_phi_mux_ack_ps
      -- 
    phi_stmt_132_phi_mux_ack_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_132_ack_0, ack => zeropad_same_CP_493_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim1_init_134_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim1_init_134_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim1_init_134_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim1_init_134_sample_start__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim1_init_134_update_start_
      -- CP-element group 46: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim1_init_134_update_start__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim1_init_134_update_completed__ps
      -- 
    zeropad_same_CP_493_elements(47) <= zeropad_same_CP_493_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim1_init_134_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => zeropad_same_CP_493_elements(46), ack => zeropad_same_CP_493_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_sample_start__ps
      -- 
    req_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(49), ack => next_input_dim1_288_135_buf_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_Update/req
      -- CP-element group 50: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_update_start_
      -- 
    req_613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(50), ack => next_input_dim1_288_135_buf_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_sample_completed_
      -- 
    ack_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim1_288_135_buf_ack_0, ack => zeropad_same_CP_493_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim1_135_update_completed_
      -- 
    ack_614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim1_288_135_buf_ack_1, ack => zeropad_same_CP_493_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: 	142 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	11 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_sample_start_
      -- 
    zeropad_same_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(142);
      gj_zeropad_same_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	133 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_update_start_
      -- 
    zeropad_same_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(133);
      gj_zeropad_same_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_sample_start__ps
      -- 
    zeropad_same_CP_493_elements(55) <= zeropad_same_CP_493_elements(11);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	13 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_update_start__ps
      -- 
    zeropad_same_CP_493_elements(57) <= zeropad_same_CP_493_elements(13);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	131 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	7 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_loopback_trigger
      -- 
    zeropad_same_CP_493_elements(59) <= zeropad_same_CP_493_elements(7);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_loopback_sample_req_ps
      -- CP-element group 60: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_loopback_sample_req
      -- 
    phi_stmt_136_loopback_sample_req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_136_loopback_sample_req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(60), ack => phi_stmt_136_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	8 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_entry_trigger
      -- 
    zeropad_same_CP_493_elements(61) <= zeropad_same_CP_493_elements(8);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_entry_sample_req_ps
      -- CP-element group 62: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_entry_sample_req
      -- 
    phi_stmt_136_entry_sample_req_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_136_entry_sample_req_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(62), ack => phi_stmt_136_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_phi_mux_ack_ps
      -- CP-element group 63: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_136_phi_mux_ack
      -- 
    phi_stmt_136_phi_mux_ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_136_ack_0, ack => zeropad_same_CP_493_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim2_init_138_sample_start__ps
      -- CP-element group 64: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim2_init_138_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim2_init_138_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim2_init_138_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim2_init_138_update_start__ps
      -- CP-element group 65: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim2_init_138_update_start_
      -- 
    -- Element group zeropad_same_CP_493_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim2_init_138_update_completed__ps
      -- 
    zeropad_same_CP_493_elements(66) <= zeropad_same_CP_493_elements(67);
    -- CP-element group 67:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	66 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_input_dim2_init_138_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => zeropad_same_CP_493_elements(65), ack => zeropad_same_CP_493_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_Sample/req
      -- CP-element group 68: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_sample_start__ps
      -- 
    req_652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(68), ack => next_input_dim2_278_139_buf_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_update_start_
      -- CP-element group 69: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_Update/req
      -- CP-element group 69: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_update_start__ps
      -- 
    req_657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(69), ack => next_input_dim2_278_139_buf_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_Sample/ack
      -- 
    ack_653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim2_278_139_buf_ack_0, ack => zeropad_same_CP_493_elements(70)); -- 
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_Update/ack
      -- CP-element group 71: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_input_dim2_139_update_completed__ps
      -- 
    ack_658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim2_278_139_buf_ack_1, ack => zeropad_same_CP_493_elements(71)); -- 
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	9 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	12 
    -- CP-element group 72: 	142 
    -- CP-element group 72: 	146 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	11 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_sample_start_
      -- 
    zeropad_same_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(142) & zeropad_same_CP_493_elements(146);
      gj_zeropad_same_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	9 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	133 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	13 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_update_start_
      -- 
    zeropad_same_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(133);
      gj_zeropad_same_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	11 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_sample_start__ps
      -- 
    zeropad_same_CP_493_elements(74) <= zeropad_same_CP_493_elements(11);
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	12 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	13 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_update_start__ps
      -- 
    zeropad_same_CP_493_elements(76) <= zeropad_same_CP_493_elements(13);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	14 
    -- CP-element group 77: 	131 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	7 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_loopback_trigger
      -- 
    zeropad_same_CP_493_elements(78) <= zeropad_same_CP_493_elements(7);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_loopback_sample_req_ps
      -- CP-element group 79: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_loopback_sample_req
      -- 
    phi_stmt_140_loopback_sample_req_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_140_loopback_sample_req_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(79), ack => phi_stmt_140_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	8 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_entry_trigger
      -- 
    zeropad_same_CP_493_elements(80) <= zeropad_same_CP_493_elements(8);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_entry_sample_req_ps
      -- CP-element group 81: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_entry_sample_req
      -- 
    phi_stmt_140_entry_sample_req_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_140_entry_sample_req_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(81), ack => phi_stmt_140_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_phi_mux_ack_ps
      -- CP-element group 82: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_140_phi_mux_ack
      -- 
    phi_stmt_140_phi_mux_ack_675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_140_ack_0, ack => zeropad_same_CP_493_elements(82)); -- 
    -- CP-element group 83:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_Sample/req
      -- CP-element group 83: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_sample_start__ps
      -- CP-element group 83: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_sample_start_
      -- 
    req_688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(83), ack => add_dest_dim0_init_118_142_buf_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_Update/req
      -- CP-element group 84: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_update_start_
      -- CP-element group 84: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_update_start__ps
      -- 
    req_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(84), ack => add_dest_dim0_init_118_142_buf_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_Sample/ack
      -- CP-element group 85: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_sample_completed__ps
      -- 
    ack_689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0_init_118_142_buf_ack_0, ack => zeropad_same_CP_493_elements(85)); -- 
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_Update/ack
      -- CP-element group 86: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim0_init_142_update_completed__ps
      -- 
    ack_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0_init_118_142_buf_ack_1, ack => zeropad_same_CP_493_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_sample_start_
      -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(87), ack => next_add_dest_dim0_272_143_buf_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_update_start_
      -- CP-element group 88: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_Update/req
      -- CP-element group 88: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_update_start__ps
      -- 
    req_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(88), ack => next_add_dest_dim0_272_143_buf_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_Sample/$exit
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim0_272_143_buf_ack_0, ack => zeropad_same_CP_493_elements(89)); -- 
    -- CP-element group 90:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_Update/ack
      -- CP-element group 90: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim0_143_update_completed__ps
      -- 
    ack_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim0_272_143_buf_ack_1, ack => zeropad_same_CP_493_elements(90)); -- 
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	9 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	12 
    -- CP-element group 91: 	142 
    -- CP-element group 91: 	146 
    -- CP-element group 91: 	150 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	11 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_sample_start_
      -- 
    zeropad_same_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(142) & zeropad_same_CP_493_elements(146) & zeropad_same_CP_493_elements(150);
      gj_zeropad_same_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	9 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	133 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	13 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_update_start_
      -- 
    zeropad_same_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad_same_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(133);
      gj_zeropad_same_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	12 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(93) is bound as output of CP function.
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: 	131 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_update_completed__ps
      -- CP-element group 94: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	7 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_loopback_trigger
      -- 
    zeropad_same_CP_493_elements(95) <= zeropad_same_CP_493_elements(7);
    -- CP-element group 96:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_loopback_sample_req
      -- CP-element group 96: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_loopback_sample_req_ps
      -- 
    phi_stmt_144_loopback_sample_req_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_144_loopback_sample_req_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(96), ack => phi_stmt_144_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	8 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_entry_trigger
      -- 
    zeropad_same_CP_493_elements(97) <= zeropad_same_CP_493_elements(8);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_entry_sample_req_ps
      -- CP-element group 98: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_entry_sample_req
      -- 
    phi_stmt_144_entry_sample_req_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_144_entry_sample_req_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(98), ack => phi_stmt_144_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_phi_mux_ack_ps
      -- CP-element group 99: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_144_phi_mux_ack
      -- 
    phi_stmt_144_phi_mux_ack_729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_144_ack_0, ack => zeropad_same_CP_493_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_Sample/req
      -- CP-element group 100: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_sample_start__ps
      -- CP-element group 100: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_Sample/$entry
      -- 
    req_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(100), ack => next_add_dest_dim1_266_146_buf_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_update_start_
      -- CP-element group 101: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_Update/req
      -- CP-element group 101: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_update_start__ps
      -- CP-element group 101: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_Update/$entry
      -- 
    req_747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(101), ack => next_add_dest_dim1_266_146_buf_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_Sample/ack
      -- CP-element group 102: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_sample_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_Sample/$exit
      -- 
    ack_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim1_266_146_buf_ack_0, ack => zeropad_same_CP_493_elements(102)); -- 
    -- CP-element group 103:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_Update/ack
      -- CP-element group 103: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_update_completed__ps
      -- CP-element group 103: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_dest_dim1_146_update_completed_
      -- 
    ack_748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim1_266_146_buf_ack_1, ack => zeropad_same_CP_493_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_Sample/req
      -- CP-element group 104: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_sample_start__ps
      -- CP-element group 104: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_sample_start_
      -- 
    req_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(104), ack => add_dest_dim1_init_121_147_buf_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_update_start__ps
      -- CP-element group 105: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_update_start_
      -- CP-element group 105: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_Update/req
      -- 
    req_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(105), ack => add_dest_dim1_init_121_147_buf_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_Sample/ack
      -- CP-element group 106: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_sample_completed_
      -- 
    ack_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1_init_121_147_buf_ack_0, ack => zeropad_same_CP_493_elements(106)); -- 
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_Update/ack
      -- CP-element group 107: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_dest_dim1_init_147_update_completed_
      -- 
    ack_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1_init_121_147_buf_ack_1, ack => zeropad_same_CP_493_elements(107)); -- 
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	9 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	12 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	11 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_sample_start_
      -- 
    zeropad_same_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(12);
      gj_zeropad_same_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	9 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	129 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	13 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_update_start_
      -- 
    zeropad_same_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(129);
      gj_zeropad_same_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	11 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_sample_start__ps
      -- 
    zeropad_same_CP_493_elements(110) <= zeropad_same_CP_493_elements(11);
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	12 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_sample_completed__ps
      -- 
    -- Element group zeropad_same_CP_493_elements(111) is bound as output of CP function.
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	13 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_update_start__ps
      -- 
    zeropad_same_CP_493_elements(112) <= zeropad_same_CP_493_elements(13);
    -- CP-element group 113:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	14 
    -- CP-element group 113: 	127 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	7 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_loopback_trigger
      -- 
    zeropad_same_CP_493_elements(114) <= zeropad_same_CP_493_elements(7);
    -- CP-element group 115:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_loopback_sample_req_ps
      -- CP-element group 115: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_loopback_sample_req
      -- 
    phi_stmt_148_loopback_sample_req_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_148_loopback_sample_req_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(115), ack => phi_stmt_148_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	8 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_entry_trigger
      -- 
    zeropad_same_CP_493_elements(116) <= zeropad_same_CP_493_elements(8);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_entry_sample_req_ps
      -- CP-element group 117: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_entry_sample_req
      -- 
    phi_stmt_148_entry_sample_req_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_148_entry_sample_req_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(117), ack => phi_stmt_148_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(117) is bound as output of CP function.
    -- CP-element group 118:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_phi_mux_ack_ps
      -- CP-element group 118: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/phi_stmt_148_phi_mux_ack
      -- 
    phi_stmt_148_phi_mux_ack_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_148_ack_0, ack => zeropad_same_CP_493_elements(118)); -- 
    -- CP-element group 119:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_src_init_150_sample_completed__ps
      -- CP-element group 119: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_src_init_150_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_src_init_150_sample_start__ps
      -- CP-element group 119: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_src_init_150_sample_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_src_init_150_update_start__ps
      -- CP-element group 120: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_src_init_150_update_start_
      -- 
    -- Element group zeropad_same_CP_493_elements(120) is bound as output of CP function.
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_src_init_150_update_completed__ps
      -- 
    zeropad_same_CP_493_elements(121) <= zeropad_same_CP_493_elements(122);
    -- CP-element group 122:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	121 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_add_src_init_150_update_completed_
      -- 
    -- Element group zeropad_same_CP_493_elements(122) is a control-delay.
    cp_element_122_delay: control_delay_element  generic map(name => " 122_delay", delay_value => 1)  port map(req => zeropad_same_CP_493_elements(120), ack => zeropad_same_CP_493_elements(122), clk => clk, reset =>reset);
    -- CP-element group 123:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_Sample/req
      -- CP-element group 123: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_sample_start__ps
      -- CP-element group 123: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_sample_start_
      -- 
    req_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(123), ack => next_add_src_253_151_buf_req_0); -- 
    -- Element group zeropad_same_CP_493_elements(123) is bound as output of CP function.
    -- CP-element group 124:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_update_start__ps
      -- CP-element group 124: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_Update/req
      -- CP-element group 124: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_update_start_
      -- 
    req_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(124), ack => next_add_src_253_151_buf_req_1); -- 
    -- Element group zeropad_same_CP_493_elements(124) is bound as output of CP function.
    -- CP-element group 125:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_sample_completed__ps
      -- CP-element group 125: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_Sample/ack
      -- CP-element group 125: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_Sample/$exit
      -- 
    ack_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_src_253_151_buf_ack_0, ack => zeropad_same_CP_493_elements(125)); -- 
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_update_completed__ps
      -- CP-element group 126: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/R_next_add_src_151_Update/ack
      -- 
    ack_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_src_253_151_buf_ack_1, ack => zeropad_same_CP_493_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	113 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_Sample/crr
      -- CP-element group 127: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_Sample/$entry
      -- 
    crr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(127), ack => call_stmt_182_call_req_0); -- 
    zeropad_same_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(113) & zeropad_same_CP_493_elements(129);
      gj_zeropad_same_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	137 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_Update/ccr
      -- CP-element group 128: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_update_start_
      -- 
    ccr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(128), ack => call_stmt_182_call_req_1); -- 
    zeropad_same_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_same_CP_493_elements(137);
      gj_zeropad_same_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	109 
    -- CP-element group 129: 	127 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_Sample/cra
      -- CP-element group 129: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_sample_completed_
      -- 
    cra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_182_call_ack_0, ack => zeropad_same_CP_493_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	135 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_Update/cca
      -- CP-element group 130: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_182_update_completed_
      -- 
    cca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_182_call_ack_1, ack => zeropad_same_CP_493_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	94 
    -- CP-element group 131: 	58 
    -- CP-element group 131: 	77 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_Sample/$entry
      -- 
    rr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(131), ack => type_cast_185_inst_req_0); -- 
    zeropad_same_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(94) & zeropad_same_CP_493_elements(58) & zeropad_same_CP_493_elements(77) & zeropad_same_CP_493_elements(133);
      gj_zeropad_same_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	137 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_update_start_
      -- CP-element group 132: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_Update/cr
      -- 
    cr_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(132), ack => type_cast_185_inst_req_1); -- 
    zeropad_same_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_same_CP_493_elements(137);
      gj_zeropad_same_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	92 
    -- CP-element group 133: 	131 
    -- CP-element group 133: 	54 
    -- CP-element group 133: 	73 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_sample_completed_
      -- 
    ra_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_0, ack => zeropad_same_CP_493_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/type_cast_185_Update/ca
      -- 
    ca_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_1, ack => zeropad_same_CP_493_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: 	130 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_Sample/crr
      -- CP-element group 135: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_sample_start_
      -- 
    crr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(135), ack => call_stmt_191_call_req_0); -- 
    zeropad_same_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(134) & zeropad_same_CP_493_elements(130) & zeropad_same_CP_493_elements(137);
      gj_zeropad_same_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_Update/ccr
      -- CP-element group 136: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_update_start_
      -- 
    ccr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(136), ack => call_stmt_191_call_req_1); -- 
    zeropad_same_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_same_CP_493_elements(138);
      gj_zeropad_same_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	132 
    -- CP-element group 137: 	135 
    -- CP-element group 137: 	128 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_Sample/cra
      -- CP-element group 137: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_sample_completed_
      -- 
    cra_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_191_call_ack_0, ack => zeropad_same_CP_493_elements(137)); -- 
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	156 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_Update/cca
      -- CP-element group 138: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/call_stmt_191_update_completed_
      -- 
    cca_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_191_call_ack_1, ack => zeropad_same_CP_493_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	9 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_Sample/req
      -- 
    req_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(139), ack => W_dim2_limit_196_delayed_1_0_197_inst_req_0); -- 
    zeropad_same_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(141);
      gj_zeropad_same_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	12 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_update_start_
      -- CP-element group 140: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_Update/req
      -- 
    req_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(140), ack => W_dim2_limit_196_delayed_1_0_197_inst_req_1); -- 
    zeropad_same_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(142);
      gj_zeropad_same_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_Sample/ack
      -- 
    ack_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dim2_limit_196_delayed_1_0_197_inst_ack_0, ack => zeropad_same_CP_493_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	10 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	91 
    -- CP-element group 142: 	15 
    -- CP-element group 142: 	34 
    -- CP-element group 142: 	140 
    -- CP-element group 142: 	53 
    -- CP-element group 142: 	72 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_199_Update/ack
      -- 
    ack_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dim2_limit_196_delayed_1_0_197_inst_ack_1, ack => zeropad_same_CP_493_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	9 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_Sample/rr
      -- 
    rr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(143), ack => SUB_u16_u16_208_inst_req_0); -- 
    zeropad_same_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(145);
      gj_zeropad_same_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	12 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_update_start_
      -- CP-element group 144: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_Update/cr
      -- 
    cr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(144), ack => SUB_u16_u16_208_inst_req_1); -- 
    zeropad_same_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(146);
      gj_zeropad_same_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_Sample/ra
      -- 
    ra_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_208_inst_ack_0, ack => zeropad_same_CP_493_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	10 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	91 
    -- CP-element group 146: 	15 
    -- CP-element group 146: 	34 
    -- CP-element group 146: 	144 
    -- CP-element group 146: 	72 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_208_Update/ca
      -- 
    ca_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_208_inst_ack_1, ack => zeropad_same_CP_493_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	9 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_Sample/req
      -- 
    req_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(147), ack => W_nid1_true4_249_delayed_1_0_254_inst_req_0); -- 
    zeropad_same_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(149);
      gj_zeropad_same_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	12 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_update_start_
      -- CP-element group 148: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_Update/req
      -- 
    req_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(148), ack => W_nid1_true4_249_delayed_1_0_254_inst_req_1); -- 
    zeropad_same_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(150);
      gj_zeropad_same_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_Sample/ack
      -- 
    ack_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_nid1_true4_249_delayed_1_0_254_inst_ack_0, ack => zeropad_same_CP_493_elements(149)); -- 
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	156 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	91 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/assign_stmt_256_Update/ack
      -- 
    ack_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_nid1_true4_249_delayed_1_0_254_inst_ack_1, ack => zeropad_same_CP_493_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	9 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_Sample/rr
      -- 
    rr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(151), ack => SUB_u16_u16_298_inst_req_0); -- 
    zeropad_same_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(9) & zeropad_same_CP_493_elements(153);
      gj_zeropad_same_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_update_start_
      -- CP-element group 152: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_Update/cr
      -- 
    cr_908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_same_CP_493_elements(152), ack => SUB_u16_u16_298_inst_req_1); -- 
    zeropad_same_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_same_CP_493_elements(154);
      gj_zeropad_same_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_Sample/ra
      -- 
    ra_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_298_inst_ack_0, ack => zeropad_same_CP_493_elements(153)); -- 
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	10 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/SUB_u16_u16_298_Update/ca
      -- 
    ca_909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_298_inst_ack_1, ack => zeropad_same_CP_493_elements(154)); -- 
    -- CP-element group 155:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	9 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	10 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group zeropad_same_CP_493_elements(155) is a control-delay.
    cp_element_155_delay: control_delay_element  generic map(name => " 155_delay", delay_value => 1)  port map(req => zeropad_same_CP_493_elements(9), ack => zeropad_same_CP_493_elements(155), clk => clk, reset =>reset);
    -- CP-element group 156:  join  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	12 
    -- CP-element group 156: 	150 
    -- CP-element group 156: 	138 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	6 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_96/do_while_stmt_126/do_while_stmt_126_loop_body/$exit
      -- 
    zeropad_same_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "zeropad_same_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_same_CP_493_elements(12) & zeropad_same_CP_493_elements(150) & zeropad_same_CP_493_elements(138);
      gj_zeropad_same_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_same_CP_493_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	5 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (2) 
      -- CP-element group 157: 	 branch_block_stmt_96/do_while_stmt_126/loop_exit/$exit
      -- CP-element group 157: 	 branch_block_stmt_96/do_while_stmt_126/loop_exit/ack
      -- 
    ack_914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_126_branch_ack_0, ack => zeropad_same_CP_493_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	5 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (2) 
      -- CP-element group 158: 	 branch_block_stmt_96/do_while_stmt_126/loop_taken/$exit
      -- CP-element group 158: 	 branch_block_stmt_96/do_while_stmt_126/loop_taken/ack
      -- 
    ack_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_126_branch_ack_1, ack => zeropad_same_CP_493_elements(158)); -- 
    -- CP-element group 159:  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	3 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	1 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_96/do_while_stmt_126/$exit
      -- 
    zeropad_same_CP_493_elements(159) <= zeropad_same_CP_493_elements(3);
    zeropad_same_do_while_stmt_126_terminator_919: loop_terminator -- 
      generic map (name => " zeropad_same_do_while_stmt_126_terminator_919", max_iterations_in_flight =>15) 
      port map(loop_body_exit => zeropad_same_CP_493_elements(6),loop_continue => zeropad_same_CP_493_elements(158),loop_terminate => zeropad_same_CP_493_elements(157),loop_back => zeropad_same_CP_493_elements(4),loop_exit => zeropad_same_CP_493_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_128_phi_seq_571_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_493_elements(23);
      zeropad_same_CP_493_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_493_elements(26);
      zeropad_same_CP_493_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_493_elements(28);
      zeropad_same_CP_493_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_493_elements(21);
      zeropad_same_CP_493_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_493_elements(32);
      zeropad_same_CP_493_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_493_elements(33);
      zeropad_same_CP_493_elements(22) <= phi_mux_reqs(1);
      phi_stmt_128_phi_seq_571 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_128_phi_seq_571") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_493_elements(17), 
          phi_sample_ack => zeropad_same_CP_493_elements(18), 
          phi_update_req => zeropad_same_CP_493_elements(19), 
          phi_update_ack => zeropad_same_CP_493_elements(20), 
          phi_mux_ack => zeropad_same_CP_493_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_132_phi_seq_615_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_493_elements(42);
      zeropad_same_CP_493_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_493_elements(45);
      zeropad_same_CP_493_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_493_elements(47);
      zeropad_same_CP_493_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_493_elements(40);
      zeropad_same_CP_493_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_493_elements(51);
      zeropad_same_CP_493_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_493_elements(52);
      zeropad_same_CP_493_elements(41) <= phi_mux_reqs(1);
      phi_stmt_132_phi_seq_615 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_132_phi_seq_615") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_493_elements(36), 
          phi_sample_ack => zeropad_same_CP_493_elements(37), 
          phi_update_req => zeropad_same_CP_493_elements(38), 
          phi_update_ack => zeropad_same_CP_493_elements(39), 
          phi_mux_ack => zeropad_same_CP_493_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_136_phi_seq_659_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_493_elements(61);
      zeropad_same_CP_493_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_493_elements(64);
      zeropad_same_CP_493_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_493_elements(66);
      zeropad_same_CP_493_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_493_elements(59);
      zeropad_same_CP_493_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_493_elements(70);
      zeropad_same_CP_493_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_493_elements(71);
      zeropad_same_CP_493_elements(60) <= phi_mux_reqs(1);
      phi_stmt_136_phi_seq_659 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_136_phi_seq_659") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_493_elements(55), 
          phi_sample_ack => zeropad_same_CP_493_elements(56), 
          phi_update_req => zeropad_same_CP_493_elements(57), 
          phi_update_ack => zeropad_same_CP_493_elements(58), 
          phi_mux_ack => zeropad_same_CP_493_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_140_phi_seq_713_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_493_elements(80);
      zeropad_same_CP_493_elements(83)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_493_elements(85);
      zeropad_same_CP_493_elements(84)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_493_elements(86);
      zeropad_same_CP_493_elements(81) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_493_elements(78);
      zeropad_same_CP_493_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_493_elements(89);
      zeropad_same_CP_493_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_493_elements(90);
      zeropad_same_CP_493_elements(79) <= phi_mux_reqs(1);
      phi_stmt_140_phi_seq_713 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_140_phi_seq_713") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_493_elements(74), 
          phi_sample_ack => zeropad_same_CP_493_elements(75), 
          phi_update_req => zeropad_same_CP_493_elements(76), 
          phi_update_ack => zeropad_same_CP_493_elements(77), 
          phi_mux_ack => zeropad_same_CP_493_elements(82), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_144_phi_seq_767_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_493_elements(95);
      zeropad_same_CP_493_elements(100)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_493_elements(102);
      zeropad_same_CP_493_elements(101)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_493_elements(103);
      zeropad_same_CP_493_elements(96) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_493_elements(97);
      zeropad_same_CP_493_elements(104)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_493_elements(106);
      zeropad_same_CP_493_elements(105)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_493_elements(107);
      zeropad_same_CP_493_elements(98) <= phi_mux_reqs(1);
      phi_stmt_144_phi_seq_767 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_144_phi_seq_767") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_493_elements(11), 
          phi_sample_ack => zeropad_same_CP_493_elements(93), 
          phi_update_req => zeropad_same_CP_493_elements(13), 
          phi_update_ack => zeropad_same_CP_493_elements(94), 
          phi_mux_ack => zeropad_same_CP_493_elements(99), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_148_phi_seq_811_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_same_CP_493_elements(116);
      zeropad_same_CP_493_elements(119)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_same_CP_493_elements(119);
      zeropad_same_CP_493_elements(120)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_same_CP_493_elements(121);
      zeropad_same_CP_493_elements(117) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_same_CP_493_elements(114);
      zeropad_same_CP_493_elements(123)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_same_CP_493_elements(125);
      zeropad_same_CP_493_elements(124)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_same_CP_493_elements(126);
      zeropad_same_CP_493_elements(115) <= phi_mux_reqs(1);
      phi_stmt_148_phi_seq_811 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_148_phi_seq_811") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_same_CP_493_elements(110), 
          phi_sample_ack => zeropad_same_CP_493_elements(111), 
          phi_update_req => zeropad_same_CP_493_elements(112), 
          phi_update_ack => zeropad_same_CP_493_elements(113), 
          phi_mux_ack => zeropad_same_CP_493_elements(118), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_523_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= zeropad_same_CP_493_elements(7);
        preds(1)  <= zeropad_same_CP_493_elements(8);
        entry_tmerge_523 : transition_merge -- 
          generic map(name => " entry_tmerge_523")
          port map (preds => preds, symbol_out => zeropad_same_CP_493_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_263_wire : std_logic_vector(15 downto 0);
    signal MUX_285_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_217_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_259_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_281_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_308_wire : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_112_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_203_203_delayed_1_0_209 : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_287_287_delayed_1_0_299 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_140 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_init_118 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_init_118_142_buffered : std_logic_vector(15 downto 0);
    signal add_dest_dim1_144 : std_logic_vector(15 downto 0);
    signal add_dest_dim1_init_121 : std_logic_vector(15 downto 0);
    signal add_dest_dim1_init_121_147_buffered : std_logic_vector(15 downto 0);
    signal add_out_177 : std_logic_vector(15 downto 0);
    signal add_src_148 : std_logic_vector(31 downto 0);
    signal add_src_init_125 : std_logic_vector(31 downto 0);
    signal cmp_dim0_220 : std_logic_vector(0 downto 0);
    signal cmp_dim1_214 : std_logic_vector(0 downto 0);
    signal cmp_dim2_204 : std_logic_vector(0 downto 0);
    signal continue_flag_310 : std_logic_vector(0 downto 0);
    signal dim0_end_304 : std_logic_vector(0 downto 0);
    signal dim2_limit_196 : std_logic_vector(15 downto 0);
    signal dim2_limit_196_delayed_1_0_199 : std_logic_vector(15 downto 0);
    signal done_191 : std_logic_vector(0 downto 0);
    signal i1_182 : std_logic_vector(63 downto 0);
    signal input_dim0_128 : std_logic_vector(15 downto 0);
    signal input_dim0_init_100 : std_logic_vector(15 downto 0);
    signal input_dim1_132 : std_logic_vector(15 downto 0);
    signal input_dim1_init_104 : std_logic_vector(15 downto 0);
    signal input_dim2_136 : std_logic_vector(15 downto 0);
    signal input_dim2_init_108 : std_logic_vector(15 downto 0);
    signal konst_113_wire_constant : std_logic_vector(15 downto 0);
    signal konst_175_wire_constant : std_logic_vector(15 downto 0);
    signal konst_194_wire_constant : std_logic_vector(15 downto 0);
    signal konst_207_wire_constant : std_logic_vector(15 downto 0);
    signal konst_223_wire_constant : std_logic_vector(15 downto 0);
    signal konst_228_wire_constant : std_logic_vector(15 downto 0);
    signal konst_233_wire_constant : std_logic_vector(15 downto 0);
    signal konst_238_wire_constant : std_logic_vector(15 downto 0);
    signal konst_243_wire_constant : std_logic_vector(15 downto 0);
    signal konst_251_wire_constant : std_logic_vector(31 downto 0);
    signal konst_276_wire_constant : std_logic_vector(15 downto 0);
    signal konst_297_wire_constant : std_logic_vector(15 downto 0);
    signal nao1_162 : std_logic_vector(15 downto 0);
    signal nao2_167 : std_logic_vector(15 downto 0);
    signal nao3_172 : std_logic_vector(15 downto 0);
    signal nao_157 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim0_272 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim0_272_143_buffered : std_logic_vector(15 downto 0);
    signal next_add_dest_dim1_266 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim1_266_146_buffered : std_logic_vector(15 downto 0);
    signal next_add_src_253 : std_logic_vector(31 downto 0);
    signal next_add_src_253_151_buffered : std_logic_vector(31 downto 0);
    signal next_input_dim0_294 : std_logic_vector(15 downto 0);
    signal next_input_dim0_294_131_buffered : std_logic_vector(15 downto 0);
    signal next_input_dim1_288 : std_logic_vector(15 downto 0);
    signal next_input_dim1_288_135_buffered : std_logic_vector(15 downto 0);
    signal next_input_dim2_278 : std_logic_vector(15 downto 0);
    signal next_input_dim2_278_139_buffered : std_logic_vector(15 downto 0);
    signal nid1_true1_245 : std_logic_vector(15 downto 0);
    signal nid1_true4_248 : std_logic_vector(15 downto 0);
    signal nid1_true4_249_delayed_1_0_256 : std_logic_vector(15 downto 0);
    signal nid1_true_240 : std_logic_vector(15 downto 0);
    signal nid2_false1_235 : std_logic_vector(15 downto 0);
    signal nid2_false_230 : std_logic_vector(15 downto 0);
    signal nid2_true_225 : std_logic_vector(15 downto 0);
    signal pad_115 : std_logic_vector(15 downto 0);
    signal type_cast_180_wire : std_logic_vector(31 downto 0);
    signal type_cast_185_185_delayed_15_0_186 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    add_src_init_125 <= "00000000000000000000000000000000";
    input_dim0_init_100 <= "0000000000000000";
    input_dim1_init_104 <= "0000000000000000";
    input_dim2_init_108 <= "0000000000000000";
    konst_113_wire_constant <= "0000000000000001";
    konst_175_wire_constant <= "0000000000000011";
    konst_194_wire_constant <= "0000000000001000";
    konst_207_wire_constant <= "0000000000000001";
    konst_223_wire_constant <= "0000000000001000";
    konst_228_wire_constant <= "0000000000000001";
    konst_233_wire_constant <= "0000000000000001";
    konst_238_wire_constant <= "0000000000000001";
    konst_243_wire_constant <= "0000000000000001";
    konst_251_wire_constant <= "00000000000000000000000000000001";
    konst_276_wire_constant <= "0000000000000000";
    konst_297_wire_constant <= "0000000000000001";
    phi_stmt_128: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim0_init_100 & next_input_dim0_294_131_buffered;
      req <= phi_stmt_128_req_0 & phi_stmt_128_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_128",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_128_ack_0,
          idata => idata,
          odata => input_dim0_128,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_128
    phi_stmt_132: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim1_init_104 & next_input_dim1_288_135_buffered;
      req <= phi_stmt_132_req_0 & phi_stmt_132_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_132",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_132_ack_0,
          idata => idata,
          odata => input_dim1_132,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_132
    phi_stmt_136: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim2_init_108 & next_input_dim2_278_139_buffered;
      req <= phi_stmt_136_req_0 & phi_stmt_136_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_136",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_136_ack_0,
          idata => idata,
          odata => input_dim2_136,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_136
    phi_stmt_140: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_dest_dim0_init_118_142_buffered & next_add_dest_dim0_272_143_buffered;
      req <= phi_stmt_140_req_0 & phi_stmt_140_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_140",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_140_ack_0,
          idata => idata,
          odata => add_dest_dim0_140,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_140
    phi_stmt_144: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_add_dest_dim1_266_146_buffered & add_dest_dim1_init_121_147_buffered;
      req <= phi_stmt_144_req_0 & phi_stmt_144_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_144",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_144_ack_0,
          idata => idata,
          odata => add_dest_dim1_144,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_144
    phi_stmt_148: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_src_init_125 & next_add_src_253_151_buffered;
      req <= phi_stmt_148_req_0 & phi_stmt_148_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_148",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_148_ack_0,
          idata => idata,
          odata => add_src_148,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_148
    -- flow-through select operator MUX_263_inst
    MUX_263_wire <= nid1_true4_249_delayed_1_0_256 when (cmp_dim1_214(0) /=  '0') else nid2_false1_235;
    -- flow-through select operator MUX_265_inst
    next_add_dest_dim1_266 <= MUX_263_wire when (NOT_u1_u1_259_wire(0) /=  '0') else add_dest_dim1_144;
    -- flow-through select operator MUX_271_inst
    next_add_dest_dim0_272 <= nid1_true1_245 when (cmp_dim0_220(0) /=  '0') else add_dest_dim0_140;
    -- flow-through select operator MUX_277_inst
    next_input_dim2_278 <= nid2_true_225 when (cmp_dim2_204(0) /=  '0') else konst_276_wire_constant;
    -- flow-through select operator MUX_285_inst
    MUX_285_wire <= pad_115 when (cmp_dim1_214(0) /=  '0') else nid2_false_230;
    -- flow-through select operator MUX_287_inst
    next_input_dim1_288 <= MUX_285_wire when (NOT_u1_u1_281_wire(0) /=  '0') else input_dim1_132;
    -- flow-through select operator MUX_293_inst
    next_input_dim0_294 <= nid1_true_240 when (cmp_dim0_220(0) /=  '0') else input_dim0_128;
    -- interlock W_add_dest_dim0_init_116_inst
    process(pad_115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := pad_115(15 downto 0);
      add_dest_dim0_init_118 <= tmp_var; -- 
    end process;
    -- interlock W_add_dest_dim1_init_119_inst
    process(pad_115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := pad_115(15 downto 0);
      add_dest_dim1_init_121 <= tmp_var; -- 
    end process;
    W_dim2_limit_196_delayed_1_0_197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_dim2_limit_196_delayed_1_0_197_inst_req_0;
      W_dim2_limit_196_delayed_1_0_197_inst_ack_0<= wack(0);
      rreq(0) <= W_dim2_limit_196_delayed_1_0_197_inst_req_1;
      W_dim2_limit_196_delayed_1_0_197_inst_ack_1<= rack(0);
      W_dim2_limit_196_delayed_1_0_197_inst : InterlockBuffer generic map ( -- 
        name => "W_dim2_limit_196_delayed_1_0_197_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => dim2_limit_196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => dim2_limit_196_delayed_1_0_199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nid1_true4_246_inst
    process(pad_115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := pad_115(15 downto 0);
      nid1_true4_248 <= tmp_var; -- 
    end process;
    W_nid1_true4_249_delayed_1_0_254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_nid1_true4_249_delayed_1_0_254_inst_req_0;
      W_nid1_true4_249_delayed_1_0_254_inst_ack_0<= wack(0);
      rreq(0) <= W_nid1_true4_249_delayed_1_0_254_inst_req_1;
      W_nid1_true4_249_delayed_1_0_254_inst_ack_1<= rack(0);
      W_nid1_true4_249_delayed_1_0_254_inst : InterlockBuffer generic map ( -- 
        name => "W_nid1_true4_249_delayed_1_0_254_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nid1_true4_248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nid1_true4_249_delayed_1_0_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim0_init_118_142_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim0_init_118_142_buf_req_0;
      add_dest_dim0_init_118_142_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim0_init_118_142_buf_req_1;
      add_dest_dim0_init_118_142_buf_ack_1<= rack(0);
      add_dest_dim0_init_118_142_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim0_init_118_142_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0_init_118,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim0_init_118_142_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim1_init_121_147_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim1_init_121_147_buf_req_0;
      add_dest_dim1_init_121_147_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim1_init_121_147_buf_req_1;
      add_dest_dim1_init_121_147_buf_ack_1<= rack(0);
      add_dest_dim1_init_121_147_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim1_init_121_147_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1_init_121,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim1_init_121_147_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_dest_dim0_272_143_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_dest_dim0_272_143_buf_req_0;
      next_add_dest_dim0_272_143_buf_ack_0<= wack(0);
      rreq(0) <= next_add_dest_dim0_272_143_buf_req_1;
      next_add_dest_dim0_272_143_buf_ack_1<= rack(0);
      next_add_dest_dim0_272_143_buf : InterlockBuffer generic map ( -- 
        name => "next_add_dest_dim0_272_143_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_dest_dim0_272,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_dest_dim0_272_143_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_dest_dim1_266_146_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_dest_dim1_266_146_buf_req_0;
      next_add_dest_dim1_266_146_buf_ack_0<= wack(0);
      rreq(0) <= next_add_dest_dim1_266_146_buf_req_1;
      next_add_dest_dim1_266_146_buf_ack_1<= rack(0);
      next_add_dest_dim1_266_146_buf : InterlockBuffer generic map ( -- 
        name => "next_add_dest_dim1_266_146_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_dest_dim1_266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_dest_dim1_266_146_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_src_253_151_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_src_253_151_buf_req_0;
      next_add_src_253_151_buf_ack_0<= wack(0);
      rreq(0) <= next_add_src_253_151_buf_req_1;
      next_add_src_253_151_buf_ack_1<= rack(0);
      next_add_src_253_151_buf : InterlockBuffer generic map ( -- 
        name => "next_add_src_253_151_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_src_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_src_253_151_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim0_294_131_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim0_294_131_buf_req_0;
      next_input_dim0_294_131_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim0_294_131_buf_req_1;
      next_input_dim0_294_131_buf_ack_1<= rack(0);
      next_input_dim0_294_131_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim0_294_131_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim0_294,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim0_294_131_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim1_288_135_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim1_288_135_buf_req_0;
      next_input_dim1_288_135_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim1_288_135_buf_req_1;
      next_input_dim1_288_135_buf_ack_1<= rack(0);
      next_input_dim1_288_135_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim1_288_135_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim1_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim1_288_135_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim2_278_139_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim2_278_139_buf_req_0;
      next_input_dim2_278_139_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim2_278_139_buf_req_1;
      next_input_dim2_278_139_buf_ack_1<= rack(0);
      next_input_dim2_278_139_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim2_278_139_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim2_278,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim2_278_139_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_180_inst
    process(add_src_148) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_src_148(31 downto 0);
      type_cast_180_wire <= tmp_var; -- 
    end process;
    type_cast_185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_185_inst_req_0;
      type_cast_185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_185_inst_req_1;
      type_cast_185_inst_ack_1<= rack(0);
      type_cast_185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_185_inst",
        buffer_size => 15,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_out_177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_185_185_delayed_15_0_186,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_126_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_310;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_126_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_126_branch_req_0,
          ack0 => do_while_stmt_126_branch_ack_0,
          ack1 => do_while_stmt_126_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_161_inst
    process(nao_157, add_dest_dim1_144) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nao_157, add_dest_dim1_144, tmp_var);
      nao1_162 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_171_inst
    process(input_dim2_136, nao2_167) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2_136, nao2_167, tmp_var);
      nao3_172 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_224_inst
    process(input_dim2_136) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2_136, konst_223_wire_constant, tmp_var);
      nid2_true_225 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_229_inst
    process(input_dim1_132) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1_132, konst_228_wire_constant, tmp_var);
      nid2_false_230 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_234_inst
    process(add_dest_dim1_144) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim1_144, konst_233_wire_constant, tmp_var);
      nid2_false1_235 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_239_inst
    process(input_dim0_128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0_128, konst_238_wire_constant, tmp_var);
      nid1_true_240 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_244_inst
    process(add_dest_dim0_140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim0_140, konst_243_wire_constant, tmp_var);
      nid1_true1_245 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_252_inst
    process(add_src_148) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_src_148, konst_251_wire_constant, tmp_var);
      next_add_src_253 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_219_inst
    process(NOT_u1_u1_217_wire, cmp_dim1_214) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_217_wire, cmp_dim1_214, tmp_var);
      cmp_dim0_220 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_213_inst
    process(input_dim1_132, SUB_u16_u16_203_203_delayed_1_0_209) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1_132, SUB_u16_u16_203_203_delayed_1_0_209, tmp_var);
      cmp_dim1_214 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_114_inst
    process(SUB_u16_u16_112_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(SUB_u16_u16_112_wire, konst_113_wire_constant, tmp_var);
      pad_115 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_176_inst
    process(nao3_172) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nao3_172, konst_175_wire_constant, tmp_var);
      add_out_177 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_156_inst
    process(out_d1_buffer, add_dest_dim0_140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d1_buffer, add_dest_dim0_140, tmp_var);
      nao_157 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_166_inst
    process(out_d2_buffer, nao1_162) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d2_buffer, nao1_162, tmp_var);
      nao2_167 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_217_inst
    process(cmp_dim2_204) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_204, tmp_var);
      NOT_u1_u1_217_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_259_inst
    process(cmp_dim2_204) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_204, tmp_var);
      NOT_u1_u1_259_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_281_inst
    process(cmp_dim2_204) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_204, tmp_var);
      NOT_u1_u1_281_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_308_inst
    process(cmp_dim0_220) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim0_220, tmp_var);
      NOT_u1_u1_308_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_309_inst
    process(dim0_end_304, NOT_u1_u1_308_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(dim0_end_304, NOT_u1_u1_308_wire, tmp_var);
      continue_flag_310 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_112_inst
    process(out_d0_buffer, inp_d0_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(out_d0_buffer, inp_d0_buffer, tmp_var);
      SUB_u16_u16_112_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_195_inst
    process(inp_d2_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(inp_d2_buffer, konst_194_wire_constant, tmp_var);
      dim2_limit_196 <= tmp_var; --
    end process;
    -- shared split operator group (21) : SUB_u16_u16_208_inst 
    ApIntSub_group_21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= inp_d1_buffer;
      SUB_u16_u16_203_203_delayed_1_0_209 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_208_inst_req_0;
      SUB_u16_u16_208_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_208_inst_req_1;
      SUB_u16_u16_208_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_21_gI: SplitGuardInterface generic map(name => "ApIntSub_group_21_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : SUB_u16_u16_298_inst 
    ApIntSub_group_22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= inp_d0_buffer;
      SUB_u16_u16_287_287_delayed_1_0_299 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_298_inst_req_0;
      SUB_u16_u16_298_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_298_inst_req_1;
      SUB_u16_u16_298_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_22_gI: SplitGuardInterface generic map(name => "ApIntSub_group_22_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- binary operator ULT_u16_u1_203_inst
    process(input_dim2_136, dim2_limit_196_delayed_1_0_199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(input_dim2_136, dim2_limit_196_delayed_1_0_199, tmp_var);
      cmp_dim2_204 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_303_inst
    process(input_dim0_128, SUB_u16_u16_287_287_delayed_1_0_299) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(input_dim0_128, SUB_u16_u16_287_287_delayed_1_0_299, tmp_var);
      dim0_end_304 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_182_call 
    readModule1_call_group_0: Block -- 
      signal data_in: std_logic_vector(39 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 15);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_182_call_req_0;
      call_stmt_182_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_182_call_req_1;
      call_stmt_182_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      readModule1_call_group_0_gI: SplitGuardInterface generic map(name => "readModule1_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= index1_buffer & type_cast_180_wire;
      i1_182 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 40,
        owidth => 40,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => readModule1_call_reqs(0),
          ackR => readModule1_call_acks(0),
          dataR => readModule1_call_data(39 downto 0),
          tagR => readModule1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => readModule1_return_acks(0), -- cross-over
          ackL => readModule1_return_reqs(0), -- cross-over
          dataL => readModule1_return_data(63 downto 0),
          tagL => readModule1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_191_call 
    writeModule1_call_group_1: Block -- 
      signal data_in: std_logic_vector(103 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 9);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_191_call_req_0;
      call_stmt_191_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_191_call_req_1;
      call_stmt_191_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeModule1_call_group_1_gI: SplitGuardInterface generic map(name => "writeModule1_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= index2_buffer & type_cast_185_185_delayed_15_0_186 & i1_182;
      done_191 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 104,
        owidth => 104,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeModule1_call_reqs(0),
          ackR => writeModule1_call_acks(0),
          dataR => writeModule1_call_data(103 downto 0),
          tagR => writeModule1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeModule1_return_acks(0), -- cross-over
          ackL => writeModule1_return_reqs(0), -- cross-over
          dataL => writeModule1_return_data(0 downto 0),
          tagL => writeModule1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad_same_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    Zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    Zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    Zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    Zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    Zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    Zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(29 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(127 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(29 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(127 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module readModule1
  component readModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(14 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readModule1
  signal readModule1_index :  std_logic_vector(7 downto 0);
  signal readModule1_address :  std_logic_vector(31 downto 0);
  signal readModule1_data :  std_logic_vector(63 downto 0);
  signal readModule1_in_args    : std_logic_vector(39 downto 0);
  signal readModule1_out_args   : std_logic_vector(63 downto 0);
  signal readModule1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal readModule1_tag_out   : std_logic_vector(1 downto 0);
  signal readModule1_start_req : std_logic;
  signal readModule1_start_ack : std_logic;
  signal readModule1_fin_req   : std_logic;
  signal readModule1_fin_ack : std_logic;
  -- caller side aggregated signals for module readModule1
  signal readModule1_call_reqs: std_logic_vector(0 downto 0);
  signal readModule1_call_acks: std_logic_vector(0 downto 0);
  signal readModule1_return_reqs: std_logic_vector(0 downto 0);
  signal readModule1_return_acks: std_logic_vector(0 downto 0);
  signal readModule1_call_data: std_logic_vector(39 downto 0);
  signal readModule1_call_tag: std_logic_vector(0 downto 0);
  signal readModule1_return_data: std_logic_vector(63 downto 0);
  signal readModule1_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- declarations related to module writeModule1
  component writeModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      done : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(14 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeModule1
  signal writeModule1_index :  std_logic_vector(7 downto 0);
  signal writeModule1_address :  std_logic_vector(31 downto 0);
  signal writeModule1_data :  std_logic_vector(63 downto 0);
  signal writeModule1_done :  std_logic_vector(0 downto 0);
  signal writeModule1_in_args    : std_logic_vector(103 downto 0);
  signal writeModule1_out_args   : std_logic_vector(0 downto 0);
  signal writeModule1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeModule1_tag_out   : std_logic_vector(1 downto 0);
  signal writeModule1_start_req : std_logic;
  signal writeModule1_start_ack : std_logic;
  signal writeModule1_fin_req   : std_logic;
  signal writeModule1_fin_ack : std_logic;
  -- caller side aggregated signals for module writeModule1
  signal writeModule1_call_reqs: std_logic_vector(0 downto 0);
  signal writeModule1_call_acks: std_logic_vector(0 downto 0);
  signal writeModule1_return_reqs: std_logic_vector(0 downto 0);
  signal writeModule1_return_acks: std_logic_vector(0 downto 0);
  signal writeModule1_call_data: std_logic_vector(103 downto 0);
  signal writeModule1_call_tag: std_logic_vector(0 downto 0);
  signal writeModule1_return_data: std_logic_vector(0 downto 0);
  signal writeModule1_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module zeropad
  component zeropad is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(14 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(14 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      Zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      Zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      zeropad_same_call_reqs : out  std_logic_vector(0 downto 0);
      zeropad_same_call_acks : in   std_logic_vector(0 downto 0);
      zeropad_same_call_data : out  std_logic_vector(111 downto 0);
      zeropad_same_call_tag  :  out  std_logic_vector(0 downto 0);
      zeropad_same_return_reqs : out  std_logic_vector(0 downto 0);
      zeropad_same_return_acks : in   std_logic_vector(0 downto 0);
      zeropad_same_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad
  signal zeropad_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad_start_req : std_logic;
  signal zeropad_start_ack : std_logic;
  signal zeropad_fin_req   : std_logic;
  signal zeropad_fin_ack : std_logic;
  -- declarations related to module zeropad_same
  component zeropad_same is -- 
    generic (tag_length : integer); 
    port ( -- 
      inp_d0 : in  std_logic_vector(15 downto 0);
      inp_d1 : in  std_logic_vector(15 downto 0);
      inp_d2 : in  std_logic_vector(15 downto 0);
      out_d0 : in  std_logic_vector(15 downto 0);
      out_d1 : in  std_logic_vector(15 downto 0);
      out_d2 : in  std_logic_vector(15 downto 0);
      index1 : in  std_logic_vector(7 downto 0);
      index2 : in  std_logic_vector(7 downto 0);
      readModule1_call_reqs : out  std_logic_vector(0 downto 0);
      readModule1_call_acks : in   std_logic_vector(0 downto 0);
      readModule1_call_data : out  std_logic_vector(39 downto 0);
      readModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      readModule1_return_reqs : out  std_logic_vector(0 downto 0);
      readModule1_return_acks : in   std_logic_vector(0 downto 0);
      readModule1_return_data : in   std_logic_vector(63 downto 0);
      readModule1_return_tag :  in   std_logic_vector(0 downto 0);
      writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_call_acks : in   std_logic_vector(0 downto 0);
      writeModule1_call_data : out  std_logic_vector(103 downto 0);
      writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_return_acks : in   std_logic_vector(0 downto 0);
      writeModule1_return_data : in   std_logic_vector(0 downto 0);
      writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad_same
  signal zeropad_same_inp_d0 :  std_logic_vector(15 downto 0);
  signal zeropad_same_inp_d1 :  std_logic_vector(15 downto 0);
  signal zeropad_same_inp_d2 :  std_logic_vector(15 downto 0);
  signal zeropad_same_out_d0 :  std_logic_vector(15 downto 0);
  signal zeropad_same_out_d1 :  std_logic_vector(15 downto 0);
  signal zeropad_same_out_d2 :  std_logic_vector(15 downto 0);
  signal zeropad_same_index1 :  std_logic_vector(7 downto 0);
  signal zeropad_same_index2 :  std_logic_vector(7 downto 0);
  signal zeropad_same_in_args    : std_logic_vector(111 downto 0);
  signal zeropad_same_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad_same_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad_same_start_req : std_logic;
  signal zeropad_same_start_ack : std_logic;
  signal zeropad_same_fin_req   : std_logic;
  signal zeropad_same_fin_ack : std_logic;
  -- caller side aggregated signals for module zeropad_same
  signal zeropad_same_call_reqs: std_logic_vector(0 downto 0);
  signal zeropad_same_call_acks: std_logic_vector(0 downto 0);
  signal zeropad_same_return_reqs: std_logic_vector(0 downto 0);
  signal zeropad_same_return_acks: std_logic_vector(0 downto 0);
  signal zeropad_same_call_data: std_logic_vector(111 downto 0);
  signal zeropad_same_call_tag: std_logic_vector(0 downto 0);
  signal zeropad_same_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Zeropad_input_pipe
  signal Zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal Zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal Zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Zeropad_output_pipe
  signal Zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal Zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal Zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module readModule1
  readModule1_index <= readModule1_in_args(39 downto 32);
  readModule1_address <= readModule1_in_args(31 downto 0);
  readModule1_out_args <= readModule1_data ;
  -- call arbiter for module readModule1
  readModule1_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 40,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => readModule1_call_reqs,
      call_acks => readModule1_call_acks,
      return_reqs => readModule1_return_reqs,
      return_acks => readModule1_return_acks,
      call_data  => readModule1_call_data,
      call_tag  => readModule1_call_tag,
      return_tag  => readModule1_return_tag,
      call_mtag => readModule1_tag_in,
      return_mtag => readModule1_tag_out,
      return_data =>readModule1_return_data,
      call_mreq => readModule1_start_req,
      call_mack => readModule1_start_ack,
      return_mreq => readModule1_fin_req,
      return_mack => readModule1_fin_ack,
      call_mdata => readModule1_in_args,
      return_mdata => readModule1_out_args,
      clk => clk, 
      reset => reset --
    ); --
  readModule1_instance:readModule1-- 
    generic map(tag_length => 2)
    port map(-- 
      index => readModule1_index,
      address => readModule1_address,
      data => readModule1_data,
      start_req => readModule1_start_req,
      start_ack => readModule1_start_ack,
      fin_req => readModule1_fin_req,
      fin_ack => readModule1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(29 downto 15),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      tag_in => readModule1_tag_in,
      tag_out => readModule1_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(0 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(0 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  -- module writeModule1
  writeModule1_index <= writeModule1_in_args(103 downto 96);
  writeModule1_address <= writeModule1_in_args(95 downto 64);
  writeModule1_data <= writeModule1_in_args(63 downto 0);
  writeModule1_out_args <= writeModule1_done ;
  -- call arbiter for module writeModule1
  writeModule1_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 104,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeModule1_call_reqs,
      call_acks => writeModule1_call_acks,
      return_reqs => writeModule1_return_reqs,
      return_acks => writeModule1_return_acks,
      call_data  => writeModule1_call_data,
      call_tag  => writeModule1_call_tag,
      return_tag  => writeModule1_return_tag,
      call_mtag => writeModule1_tag_in,
      return_mtag => writeModule1_tag_out,
      return_data =>writeModule1_return_data,
      call_mreq => writeModule1_start_req,
      call_mack => writeModule1_start_ack,
      return_mreq => writeModule1_fin_req,
      return_mack => writeModule1_fin_ack,
      call_mdata => writeModule1_in_args,
      return_mdata => writeModule1_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeModule1_instance:writeModule1-- 
    generic map(tag_length => 2)
    port map(-- 
      index => writeModule1_index,
      address => writeModule1_address,
      data => writeModule1_data,
      done => writeModule1_done,
      start_req => writeModule1_start_req,
      start_ack => writeModule1_start_ack,
      fin_req => writeModule1_fin_req,
      fin_ack => writeModule1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(29 downto 15),
      memory_space_0_sr_data => memory_space_0_sr_data(127 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(39 downto 20),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      tag_in => writeModule1_tag_in,
      tag_out => writeModule1_tag_out-- 
    ); -- 
  -- module zeropad
  zeropad_instance:zeropad-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad_start_req,
      start_ack => zeropad_start_ack,
      fin_req => zeropad_fin_req,
      fin_ack => zeropad_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(14 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(14 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      Zeropad_input_pipe_pipe_read_req => Zeropad_input_pipe_pipe_read_req(0 downto 0),
      Zeropad_input_pipe_pipe_read_ack => Zeropad_input_pipe_pipe_read_ack(0 downto 0),
      Zeropad_input_pipe_pipe_read_data => Zeropad_input_pipe_pipe_read_data(7 downto 0),
      Zeropad_output_pipe_pipe_write_req => Zeropad_output_pipe_pipe_write_req(0 downto 0),
      Zeropad_output_pipe_pipe_write_ack => Zeropad_output_pipe_pipe_write_ack(0 downto 0),
      Zeropad_output_pipe_pipe_write_data => Zeropad_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      zeropad_same_call_reqs => zeropad_same_call_reqs(0 downto 0),
      zeropad_same_call_acks => zeropad_same_call_acks(0 downto 0),
      zeropad_same_call_data => zeropad_same_call_data(111 downto 0),
      zeropad_same_call_tag => zeropad_same_call_tag(0 downto 0),
      zeropad_same_return_reqs => zeropad_same_return_reqs(0 downto 0),
      zeropad_same_return_acks => zeropad_same_return_acks(0 downto 0),
      zeropad_same_return_tag => zeropad_same_return_tag(0 downto 0),
      tag_in => zeropad_tag_in,
      tag_out => zeropad_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad_tag_in <= (others => '0');
  zeropad_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad_start_req, start_ack => zeropad_start_ack,  fin_req => zeropad_fin_req,  fin_ack => zeropad_fin_ack);
  -- module zeropad_same
  zeropad_same_inp_d0 <= zeropad_same_in_args(111 downto 96);
  zeropad_same_inp_d1 <= zeropad_same_in_args(95 downto 80);
  zeropad_same_inp_d2 <= zeropad_same_in_args(79 downto 64);
  zeropad_same_out_d0 <= zeropad_same_in_args(63 downto 48);
  zeropad_same_out_d1 <= zeropad_same_in_args(47 downto 32);
  zeropad_same_out_d2 <= zeropad_same_in_args(31 downto 16);
  zeropad_same_index1 <= zeropad_same_in_args(15 downto 8);
  zeropad_same_index2 <= zeropad_same_in_args(7 downto 0);
  -- call arbiter for module zeropad_same
  zeropad_same_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 112,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => zeropad_same_call_reqs,
      call_acks => zeropad_same_call_acks,
      return_reqs => zeropad_same_return_reqs,
      return_acks => zeropad_same_return_acks,
      call_data  => zeropad_same_call_data,
      call_tag  => zeropad_same_call_tag,
      return_tag  => zeropad_same_return_tag,
      call_mtag => zeropad_same_tag_in,
      return_mtag => zeropad_same_tag_out,
      call_mreq => zeropad_same_start_req,
      call_mack => zeropad_same_start_ack,
      return_mreq => zeropad_same_fin_req,
      return_mack => zeropad_same_fin_ack,
      call_mdata => zeropad_same_in_args,
      clk => clk, 
      reset => reset --
    ); --
  zeropad_same_instance:zeropad_same-- 
    generic map(tag_length => 2)
    port map(-- 
      inp_d0 => zeropad_same_inp_d0,
      inp_d1 => zeropad_same_inp_d1,
      inp_d2 => zeropad_same_inp_d2,
      out_d0 => zeropad_same_out_d0,
      out_d1 => zeropad_same_out_d1,
      out_d2 => zeropad_same_out_d2,
      index1 => zeropad_same_index1,
      index2 => zeropad_same_index2,
      start_req => zeropad_same_start_req,
      start_ack => zeropad_same_start_ack,
      fin_req => zeropad_same_fin_req,
      fin_ack => zeropad_same_fin_ack,
      clk => clk,
      reset => reset,
      readModule1_call_reqs => readModule1_call_reqs(0 downto 0),
      readModule1_call_acks => readModule1_call_acks(0 downto 0),
      readModule1_call_data => readModule1_call_data(39 downto 0),
      readModule1_call_tag => readModule1_call_tag(0 downto 0),
      readModule1_return_reqs => readModule1_return_reqs(0 downto 0),
      readModule1_return_acks => readModule1_return_acks(0 downto 0),
      readModule1_return_data => readModule1_return_data(63 downto 0),
      readModule1_return_tag => readModule1_return_tag(0 downto 0),
      writeModule1_call_reqs => writeModule1_call_reqs(0 downto 0),
      writeModule1_call_acks => writeModule1_call_acks(0 downto 0),
      writeModule1_call_data => writeModule1_call_data(103 downto 0),
      writeModule1_call_tag => writeModule1_call_tag(0 downto 0),
      writeModule1_return_reqs => writeModule1_return_reqs(0 downto 0),
      writeModule1_return_acks => writeModule1_return_acks(0 downto 0),
      writeModule1_return_data => writeModule1_return_data(0 downto 0),
      writeModule1_return_tag => writeModule1_return_tag(0 downto 0),
      tag_in => zeropad_same_tag_in,
      tag_out => zeropad_same_tag_out-- 
    ); -- 
  Zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Zeropad_input_pipe_pipe_read_req,
      read_ack => Zeropad_input_pipe_pipe_read_ack,
      read_data => Zeropad_input_pipe_pipe_read_data,
      write_req => Zeropad_input_pipe_pipe_write_req,
      write_ack => Zeropad_input_pipe_pipe_write_ack,
      write_data => Zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Zeropad_output_pipe_pipe_read_req,
      read_ack => Zeropad_output_pipe_pipe_read_ack,
      read_data => Zeropad_output_pipe_pipe_read_data,
      write_req => Zeropad_output_pipe_pipe_write_req,
      write_ack => Zeropad_output_pipe_pipe_write_ack,
      write_data => Zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 2,
      addr_width => 15,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 15,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
