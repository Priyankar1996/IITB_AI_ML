-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    row_in : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe4_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 48)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal row_in_buffer :  std_logic_vector(15 downto 0);
  signal row_in_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal W_send3_1_280_delayed_14_0_286_inst_req_1 : boolean;
  signal slice_504_inst_req_0 : boolean;
  signal slice_504_inst_req_1 : boolean;
  signal W_send1_1_272_delayed_14_0_272_inst_req_1 : boolean;
  signal WPIPE_input_pipe3_634_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_283_inst_req_0 : boolean;
  signal W_send2_3_596_delayed_14_0_623_inst_ack_1 : boolean;
  signal slice_676_inst_req_1 : boolean;
  signal n_start3_512_120_buf_ack_0 : boolean;
  signal W_send4_1_284_delayed_14_0_293_inst_req_1 : boolean;
  signal W_send4_1_284_delayed_14_0_293_inst_ack_1 : boolean;
  signal W_send4_1_284_delayed_14_0_293_inst_req_0 : boolean;
  signal W_send4_1_284_delayed_14_0_293_inst_ack_0 : boolean;
  signal W_send3_1_280_delayed_14_0_286_inst_ack_1 : boolean;
  signal n_start4_684_125_buf_ack_1 : boolean;
  signal phi_stmt_44_req_0 : boolean;
  signal n_start3_512_120_buf_req_0 : boolean;
  signal do_while_stmt_42_branch_req_0 : boolean;
  signal slice_492_inst_req_1 : boolean;
  signal slice_159_inst_ack_1 : boolean;
  signal phi_stmt_44_req_1 : boolean;
  signal W_send3_1_280_delayed_14_0_286_inst_ack_0 : boolean;
  signal slice_155_inst_ack_1 : boolean;
  signal phi_stmt_44_ack_0 : boolean;
  signal slice_155_inst_req_1 : boolean;
  signal n_address1_210_48_buf_req_0 : boolean;
  signal n_address1_210_48_buf_ack_0 : boolean;
  signal n_address1_210_48_buf_req_1 : boolean;
  signal n_address1_210_48_buf_ack_1 : boolean;
  signal n_start4_684_125_buf_ack_0 : boolean;
  signal n_start4_684_125_buf_req_0 : boolean;
  signal slice_159_inst_req_1 : boolean;
  signal slice_147_inst_ack_1 : boolean;
  signal slice_664_inst_req_1 : boolean;
  signal phi_stmt_49_req_0 : boolean;
  signal slice_147_inst_req_1 : boolean;
  signal phi_stmt_49_req_1 : boolean;
  signal slice_147_inst_ack_0 : boolean;
  signal W_send3_1_280_delayed_14_0_286_inst_req_0 : boolean;
  signal slice_155_inst_ack_0 : boolean;
  signal phi_stmt_49_ack_0 : boolean;
  signal W_send1_1_272_delayed_14_0_272_inst_ack_0 : boolean;
  signal W_send4_3_604_delayed_14_0_637_inst_req_1 : boolean;
  signal n_address2_382_51_buf_req_0 : boolean;
  signal n_address2_382_51_buf_ack_0 : boolean;
  signal slice_147_inst_req_0 : boolean;
  signal n_address2_382_51_buf_req_1 : boolean;
  signal n_address2_382_51_buf_ack_1 : boolean;
  signal slice_155_inst_req_0 : boolean;
  signal phi_stmt_66_req_0 : boolean;
  signal phi_stmt_66_ack_0 : boolean;
  signal W_send1_3_592_delayed_14_0_616_inst_ack_0 : boolean;
  signal type_cast_53_inst_req_0 : boolean;
  signal type_cast_53_inst_ack_0 : boolean;
  signal type_cast_53_inst_req_1 : boolean;
  signal array_obj_ref_655_index_offset_req_1 : boolean;
  signal type_cast_53_inst_ack_1 : boolean;
  signal WPIPE_input_pipe3_634_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_276_inst_ack_1 : boolean;
  signal slice_672_inst_ack_0 : boolean;
  signal n_start4_684_125_buf_req_1 : boolean;
  signal WPIPE_input_pipe1_276_inst_req_1 : boolean;
  signal phi_stmt_54_req_0 : boolean;
  signal WPIPE_input_pipe1_290_inst_ack_0 : boolean;
  signal phi_stmt_54_req_1 : boolean;
  signal phi_stmt_54_ack_0 : boolean;
  signal W_send1_1_272_delayed_14_0_272_inst_req_0 : boolean;
  signal addr_of_139_final_reg_ack_1 : boolean;
  signal addr_of_139_final_reg_req_1 : boolean;
  signal n_address3_554_56_buf_req_0 : boolean;
  signal n_address3_554_56_buf_ack_0 : boolean;
  signal n_address3_554_56_buf_req_1 : boolean;
  signal n_address3_554_56_buf_ack_1 : boolean;
  signal WPIPE_input_pipe1_276_inst_ack_0 : boolean;
  signal addr_of_139_final_reg_ack_0 : boolean;
  signal addr_of_139_final_reg_req_0 : boolean;
  signal type_cast_58_inst_req_0 : boolean;
  signal type_cast_58_inst_ack_0 : boolean;
  signal type_cast_58_inst_req_1 : boolean;
  signal type_cast_58_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_276_inst_req_0 : boolean;
  signal slice_159_inst_ack_0 : boolean;
  signal slice_159_inst_req_0 : boolean;
  signal phi_stmt_59_req_1 : boolean;
  signal WPIPE_input_pipe1_290_inst_req_0 : boolean;
  signal phi_stmt_59_req_0 : boolean;
  signal W_send1_3_592_delayed_14_0_616_inst_req_0 : boolean;
  signal phi_stmt_59_ack_0 : boolean;
  signal ptr_deref_488_load_0_req_0 : boolean;
  signal ptr_deref_488_load_0_ack_0 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal array_obj_ref_655_index_offset_ack_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal slice_668_inst_ack_1 : boolean;
  signal n_address4_726_65_buf_req_0 : boolean;
  signal n_address4_726_65_buf_ack_0 : boolean;
  signal n_address4_726_65_buf_req_1 : boolean;
  signal n_address4_726_65_buf_ack_1 : boolean;
  signal slice_668_inst_req_1 : boolean;
  signal slice_676_inst_ack_1 : boolean;
  signal W_send4_3_604_delayed_14_0_637_inst_ack_1 : boolean;
  signal phi_stmt_66_req_1 : boolean;
  signal phi_stmt_121_req_1 : boolean;
  signal n_row2_365_95_buf_req_0 : boolean;
  signal n_row2_365_95_buf_ack_0 : boolean;
  signal phi_stmt_116_req_1 : boolean;
  signal n_row2_365_95_buf_req_1 : boolean;
  signal n_row2_365_95_buf_ack_1 : boolean;
  signal type_cast_69_inst_req_0 : boolean;
  signal type_cast_69_inst_ack_0 : boolean;
  signal WPIPE_input_pipe3_627_inst_req_1 : boolean;
  signal type_cast_69_inst_req_1 : boolean;
  signal type_cast_69_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_283_inst_ack_1 : boolean;
  signal array_obj_ref_138_index_offset_ack_1 : boolean;
  signal array_obj_ref_138_index_offset_req_1 : boolean;
  signal n_mycounter1_185_70_buf_req_0 : boolean;
  signal n_mycounter1_185_70_buf_ack_0 : boolean;
  signal slice_504_inst_ack_1 : boolean;
  signal n_mycounter1_185_70_buf_req_1 : boolean;
  signal n_mycounter1_185_70_buf_ack_1 : boolean;
  signal WPIPE_input_pipe1_283_inst_req_1 : boolean;
  signal array_obj_ref_655_index_offset_req_0 : boolean;
  signal phi_stmt_71_req_1 : boolean;
  signal phi_stmt_71_req_0 : boolean;
  signal ptr_deref_143_load_0_ack_1 : boolean;
  signal W_send2_1_276_delayed_14_0_279_inst_ack_1 : boolean;
  signal array_obj_ref_655_index_offset_ack_0 : boolean;
  signal phi_stmt_71_ack_0 : boolean;
  signal array_obj_ref_138_index_offset_ack_0 : boolean;
  signal array_obj_ref_138_index_offset_req_0 : boolean;
  signal type_cast_74_inst_req_0 : boolean;
  signal type_cast_74_inst_ack_0 : boolean;
  signal ptr_deref_143_load_0_req_1 : boolean;
  signal type_cast_74_inst_req_1 : boolean;
  signal type_cast_74_inst_ack_1 : boolean;
  signal slice_504_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_290_inst_ack_1 : boolean;
  signal n_mycounter2_357_75_buf_req_0 : boolean;
  signal n_mycounter2_357_75_buf_ack_0 : boolean;
  signal W_send2_1_276_delayed_14_0_279_inst_req_1 : boolean;
  signal n_mycounter2_357_75_buf_req_1 : boolean;
  signal n_mycounter2_357_75_buf_ack_1 : boolean;
  signal WPIPE_input_pipe4_792_inst_ack_0 : boolean;
  signal n_start3_512_120_buf_ack_1 : boolean;
  signal phi_stmt_76_req_1 : boolean;
  signal phi_stmt_76_req_0 : boolean;
  signal phi_stmt_76_ack_0 : boolean;
  signal type_cast_79_inst_req_0 : boolean;
  signal type_cast_79_inst_ack_0 : boolean;
  signal type_cast_79_inst_req_1 : boolean;
  signal type_cast_79_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_290_inst_req_1 : boolean;
  signal slice_672_inst_req_0 : boolean;
  signal n_mycounter3_529_80_buf_req_0 : boolean;
  signal n_mycounter3_529_80_buf_ack_0 : boolean;
  signal n_mycounter3_529_80_buf_req_1 : boolean;
  signal n_mycounter3_529_80_buf_ack_1 : boolean;
  signal n_start3_512_120_buf_req_1 : boolean;
  signal WPIPE_input_pipe1_283_inst_ack_0 : boolean;
  signal ptr_deref_143_load_0_ack_0 : boolean;
  signal ptr_deref_143_load_0_req_0 : boolean;
  signal slice_664_inst_ack_1 : boolean;
  signal W_send1_1_272_delayed_14_0_272_inst_ack_1 : boolean;
  signal phi_stmt_81_req_1 : boolean;
  signal WPIPE_input_pipe4_792_inst_req_0 : boolean;
  signal phi_stmt_81_req_0 : boolean;
  signal W_send2_1_276_delayed_14_0_279_inst_ack_0 : boolean;
  signal W_send4_3_604_delayed_14_0_637_inst_req_0 : boolean;
  signal phi_stmt_81_ack_0 : boolean;
  signal slice_151_inst_ack_1 : boolean;
  signal W_send1_3_592_delayed_14_0_616_inst_req_1 : boolean;
  signal type_cast_84_inst_req_0 : boolean;
  signal slice_492_inst_ack_1 : boolean;
  signal type_cast_84_inst_ack_0 : boolean;
  signal type_cast_84_inst_req_1 : boolean;
  signal type_cast_84_inst_ack_1 : boolean;
  signal W_send1_4_752_delayed_14_0_788_inst_ack_1 : boolean;
  signal W_send4_3_604_delayed_14_0_637_inst_ack_0 : boolean;
  signal W_send1_3_592_delayed_14_0_616_inst_ack_1 : boolean;
  signal n_mycounter4_701_85_buf_req_0 : boolean;
  signal n_mycounter4_701_85_buf_ack_0 : boolean;
  signal W_send2_1_276_delayed_14_0_279_inst_req_0 : boolean;
  signal n_mycounter4_701_85_buf_req_1 : boolean;
  signal n_mycounter4_701_85_buf_ack_1 : boolean;
  signal phi_stmt_116_ack_0 : boolean;
  signal phi_stmt_86_req_0 : boolean;
  signal slice_151_inst_req_1 : boolean;
  signal phi_stmt_86_req_1 : boolean;
  signal phi_stmt_86_ack_0 : boolean;
  signal phi_stmt_121_ack_0 : boolean;
  signal n_row1_193_88_buf_req_0 : boolean;
  signal n_row1_193_88_buf_ack_0 : boolean;
  signal phi_stmt_116_req_0 : boolean;
  signal n_row1_193_88_buf_req_1 : boolean;
  signal n_row1_193_88_buf_ack_1 : boolean;
  signal slice_151_inst_ack_0 : boolean;
  signal phi_stmt_121_req_0 : boolean;
  signal slice_151_inst_req_0 : boolean;
  signal slice_492_inst_req_0 : boolean;
  signal phi_stmt_91_req_1 : boolean;
  signal phi_stmt_91_req_0 : boolean;
  signal ptr_deref_488_load_0_req_1 : boolean;
  signal phi_stmt_91_ack_0 : boolean;
  signal ptr_deref_488_load_0_ack_1 : boolean;
  signal WPIPE_input_pipe3_627_inst_req_0 : boolean;
  signal phi_stmt_96_req_1 : boolean;
  signal ptr_deref_660_load_0_req_0 : boolean;
  signal phi_stmt_96_req_0 : boolean;
  signal WPIPE_input_pipe3_641_inst_req_0 : boolean;
  signal phi_stmt_96_ack_0 : boolean;
  signal WPIPE_input_pipe3_641_inst_ack_0 : boolean;
  signal n_row3_537_100_buf_req_0 : boolean;
  signal n_row3_537_100_buf_ack_0 : boolean;
  signal n_row3_537_100_buf_req_1 : boolean;
  signal n_row3_537_100_buf_ack_1 : boolean;
  signal WPIPE_input_pipe3_620_inst_req_0 : boolean;
  signal WPIPE_input_pipe3_627_inst_ack_0 : boolean;
  signal WPIPE_input_pipe3_620_inst_ack_0 : boolean;
  signal ptr_deref_660_load_0_ack_0 : boolean;
  signal phi_stmt_101_req_1 : boolean;
  signal phi_stmt_101_req_0 : boolean;
  signal phi_stmt_101_ack_0 : boolean;
  signal WPIPE_input_pipe3_641_inst_req_1 : boolean;
  signal WPIPE_input_pipe3_641_inst_ack_1 : boolean;
  signal WPIPE_input_pipe3_620_inst_req_1 : boolean;
  signal WPIPE_input_pipe3_620_inst_ack_1 : boolean;
  signal n_row4_709_105_buf_req_0 : boolean;
  signal n_row4_709_105_buf_ack_0 : boolean;
  signal n_row4_709_105_buf_req_1 : boolean;
  signal n_row4_709_105_buf_ack_1 : boolean;
  signal phi_stmt_106_req_1 : boolean;
  signal phi_stmt_106_req_0 : boolean;
  signal phi_stmt_106_ack_0 : boolean;
  signal n_start1_168_110_buf_req_0 : boolean;
  signal n_start1_168_110_buf_ack_0 : boolean;
  signal n_start1_168_110_buf_req_1 : boolean;
  signal n_start1_168_110_buf_ack_1 : boolean;
  signal phi_stmt_111_req_1 : boolean;
  signal phi_stmt_111_req_0 : boolean;
  signal phi_stmt_111_ack_0 : boolean;
  signal n_start2_340_115_buf_req_0 : boolean;
  signal n_start2_340_115_buf_ack_0 : boolean;
  signal n_start2_340_115_buf_req_1 : boolean;
  signal n_start2_340_115_buf_ack_1 : boolean;
  signal W_send1_4_752_delayed_14_0_788_inst_ack_0 : boolean;
  signal W_send2_4_756_delayed_14_0_795_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_297_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_297_inst_ack_0 : boolean;
  signal slice_500_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_297_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_297_inst_ack_1 : boolean;
  signal W_send2_3_596_delayed_14_0_623_inst_req_1 : boolean;
  signal addr_of_656_final_reg_ack_1 : boolean;
  signal addr_of_656_final_reg_req_1 : boolean;
  signal WPIPE_input_pipe3_634_inst_ack_0 : boolean;
  signal WPIPE_input_pipe3_634_inst_req_0 : boolean;
  signal array_obj_ref_311_index_offset_req_0 : boolean;
  signal array_obj_ref_311_index_offset_ack_0 : boolean;
  signal slice_500_inst_req_1 : boolean;
  signal array_obj_ref_311_index_offset_req_1 : boolean;
  signal array_obj_ref_311_index_offset_ack_1 : boolean;
  signal slice_664_inst_ack_0 : boolean;
  signal addr_of_312_final_reg_req_0 : boolean;
  signal addr_of_312_final_reg_ack_0 : boolean;
  signal addr_of_312_final_reg_req_1 : boolean;
  signal addr_of_312_final_reg_ack_1 : boolean;
  signal W_send1_4_752_delayed_14_0_788_inst_req_1 : boolean;
  signal slice_668_inst_ack_0 : boolean;
  signal W_send1_4_752_delayed_14_0_788_inst_req_0 : boolean;
  signal addr_of_656_final_reg_ack_0 : boolean;
  signal addr_of_656_final_reg_req_0 : boolean;
  signal W_send2_3_596_delayed_14_0_623_inst_ack_0 : boolean;
  signal ptr_deref_316_load_0_req_0 : boolean;
  signal ptr_deref_316_load_0_ack_0 : boolean;
  signal slice_492_inst_ack_0 : boolean;
  signal W_send2_3_596_delayed_14_0_623_inst_req_0 : boolean;
  signal ptr_deref_316_load_0_req_1 : boolean;
  signal ptr_deref_316_load_0_ack_1 : boolean;
  signal W_send3_3_600_delayed_14_0_630_inst_ack_1 : boolean;
  signal slice_668_inst_req_0 : boolean;
  signal slice_664_inst_req_0 : boolean;
  signal W_send3_3_600_delayed_14_0_630_inst_req_1 : boolean;
  signal slice_320_inst_req_0 : boolean;
  signal slice_320_inst_ack_0 : boolean;
  signal slice_320_inst_req_1 : boolean;
  signal slice_320_inst_ack_1 : boolean;
  signal slice_500_inst_ack_0 : boolean;
  signal slice_324_inst_req_0 : boolean;
  signal slice_324_inst_ack_0 : boolean;
  signal slice_324_inst_req_1 : boolean;
  signal slice_324_inst_ack_1 : boolean;
  signal slice_500_inst_req_0 : boolean;
  signal slice_328_inst_req_0 : boolean;
  signal slice_328_inst_ack_0 : boolean;
  signal slice_328_inst_req_1 : boolean;
  signal slice_328_inst_ack_1 : boolean;
  signal slice_332_inst_req_0 : boolean;
  signal slice_332_inst_ack_0 : boolean;
  signal slice_332_inst_req_1 : boolean;
  signal slice_332_inst_ack_1 : boolean;
  signal W_send1_2_432_delayed_14_0_444_inst_req_0 : boolean;
  signal W_send1_2_432_delayed_14_0_444_inst_ack_0 : boolean;
  signal W_send1_2_432_delayed_14_0_444_inst_req_1 : boolean;
  signal W_send1_2_432_delayed_14_0_444_inst_ack_1 : boolean;
  signal WPIPE_input_pipe4_792_inst_ack_1 : boolean;
  signal W_send2_4_756_delayed_14_0_795_inst_ack_1 : boolean;
  signal ptr_deref_660_load_0_ack_1 : boolean;
  signal WPIPE_input_pipe2_448_inst_req_0 : boolean;
  signal WPIPE_input_pipe2_448_inst_ack_0 : boolean;
  signal WPIPE_input_pipe2_448_inst_req_1 : boolean;
  signal WPIPE_input_pipe2_448_inst_ack_1 : boolean;
  signal ptr_deref_660_load_0_req_1 : boolean;
  signal W_send2_2_436_delayed_14_0_451_inst_req_0 : boolean;
  signal W_send2_2_436_delayed_14_0_451_inst_ack_0 : boolean;
  signal W_send2_2_436_delayed_14_0_451_inst_req_1 : boolean;
  signal W_send2_2_436_delayed_14_0_451_inst_ack_1 : boolean;
  signal WPIPE_input_pipe4_792_inst_req_1 : boolean;
  signal W_send2_4_756_delayed_14_0_795_inst_req_0 : boolean;
  signal WPIPE_input_pipe2_455_inst_req_0 : boolean;
  signal WPIPE_input_pipe2_455_inst_ack_0 : boolean;
  signal WPIPE_input_pipe2_455_inst_req_1 : boolean;
  signal WPIPE_input_pipe2_455_inst_ack_1 : boolean;
  signal W_send3_3_600_delayed_14_0_630_inst_ack_0 : boolean;
  signal W_send3_2_440_delayed_14_0_458_inst_req_0 : boolean;
  signal W_send3_2_440_delayed_14_0_458_inst_ack_0 : boolean;
  signal W_send3_2_440_delayed_14_0_458_inst_req_1 : boolean;
  signal W_send3_2_440_delayed_14_0_458_inst_ack_1 : boolean;
  signal slice_676_inst_ack_0 : boolean;
  signal slice_676_inst_req_0 : boolean;
  signal W_send2_4_756_delayed_14_0_795_inst_ack_0 : boolean;
  signal slice_496_inst_ack_1 : boolean;
  signal slice_672_inst_ack_1 : boolean;
  signal WPIPE_input_pipe2_462_inst_req_0 : boolean;
  signal WPIPE_input_pipe2_462_inst_ack_0 : boolean;
  signal slice_496_inst_req_1 : boolean;
  signal WPIPE_input_pipe2_462_inst_req_1 : boolean;
  signal WPIPE_input_pipe2_462_inst_ack_1 : boolean;
  signal W_send3_3_600_delayed_14_0_630_inst_req_0 : boolean;
  signal W_send4_2_444_delayed_14_0_465_inst_req_0 : boolean;
  signal W_send4_2_444_delayed_14_0_465_inst_ack_0 : boolean;
  signal W_send4_2_444_delayed_14_0_465_inst_req_1 : boolean;
  signal W_send4_2_444_delayed_14_0_465_inst_ack_1 : boolean;
  signal slice_672_inst_req_1 : boolean;
  signal slice_496_inst_ack_0 : boolean;
  signal WPIPE_input_pipe2_469_inst_req_0 : boolean;
  signal WPIPE_input_pipe2_469_inst_ack_0 : boolean;
  signal slice_496_inst_req_0 : boolean;
  signal WPIPE_input_pipe2_469_inst_req_1 : boolean;
  signal WPIPE_input_pipe2_469_inst_ack_1 : boolean;
  signal WPIPE_input_pipe3_627_inst_ack_1 : boolean;
  signal array_obj_ref_483_index_offset_req_0 : boolean;
  signal array_obj_ref_483_index_offset_ack_0 : boolean;
  signal array_obj_ref_483_index_offset_req_1 : boolean;
  signal array_obj_ref_483_index_offset_ack_1 : boolean;
  signal addr_of_484_final_reg_req_0 : boolean;
  signal addr_of_484_final_reg_ack_0 : boolean;
  signal addr_of_484_final_reg_req_1 : boolean;
  signal addr_of_484_final_reg_ack_1 : boolean;
  signal WPIPE_input_pipe4_799_inst_req_0 : boolean;
  signal WPIPE_input_pipe4_799_inst_ack_0 : boolean;
  signal WPIPE_input_pipe4_799_inst_req_1 : boolean;
  signal WPIPE_input_pipe4_799_inst_ack_1 : boolean;
  signal W_send3_4_760_delayed_14_0_802_inst_req_0 : boolean;
  signal W_send3_4_760_delayed_14_0_802_inst_ack_0 : boolean;
  signal W_send3_4_760_delayed_14_0_802_inst_req_1 : boolean;
  signal W_send3_4_760_delayed_14_0_802_inst_ack_1 : boolean;
  signal WPIPE_input_pipe4_806_inst_req_0 : boolean;
  signal WPIPE_input_pipe4_806_inst_ack_0 : boolean;
  signal WPIPE_input_pipe4_806_inst_req_1 : boolean;
  signal WPIPE_input_pipe4_806_inst_ack_1 : boolean;
  signal W_send4_4_764_delayed_14_0_809_inst_req_0 : boolean;
  signal W_send4_4_764_delayed_14_0_809_inst_ack_0 : boolean;
  signal W_send4_4_764_delayed_14_0_809_inst_req_1 : boolean;
  signal W_send4_4_764_delayed_14_0_809_inst_ack_1 : boolean;
  signal WPIPE_input_pipe4_813_inst_req_0 : boolean;
  signal WPIPE_input_pipe4_813_inst_ack_0 : boolean;
  signal WPIPE_input_pipe4_813_inst_req_1 : boolean;
  signal WPIPE_input_pipe4_813_inst_ack_1 : boolean;
  signal do_while_stmt_42_branch_ack_0 : boolean;
  signal do_while_stmt_42_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 48) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= row_in;
  row_in_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= ct;
  ct_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(tag_length + 47 downto 48) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 47 downto 48);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(555 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_41__exit__
      -- CP-element group 0: 	 branch_block_stmt_29/do_while_stmt_42__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_41/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_41/$exit
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_29/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/branch_block_stmt_29__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_41__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	555 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_29/do_while_stmt_42__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_29/$exit
      -- CP-element group 1: 	 branch_block_stmt_29/branch_block_stmt_29__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(555);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_29/do_while_stmt_42/$entry
      -- CP-element group 2: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	555 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_29/do_while_stmt_42/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	553 
    -- CP-element group 5: 	554 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_29/do_while_stmt_42/condition_done
      -- CP-element group 5: 	 branch_block_stmt_29/do_while_stmt_42/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_29/do_while_stmt_42/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	552 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_29/do_while_stmt_42/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(552);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	280 
    -- CP-element group 7: 	145 
    -- CP-element group 7: 	187 
    -- CP-element group 7: 	166 
    -- CP-element group 7: 	299 
    -- CP-element group 7: 	318 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	61 
    -- CP-element group 7: 	82 
    -- CP-element group 7: 	206 
    -- CP-element group 7: 	225 
    -- CP-element group 7: 	244 
    -- CP-element group 7: 	263 
    -- CP-element group 7: 	103 
    -- CP-element group 7: 	124 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	282 
    -- CP-element group 8: 	147 
    -- CP-element group 8: 	189 
    -- CP-element group 8: 	168 
    -- CP-element group 8: 	301 
    -- CP-element group 8: 	320 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	63 
    -- CP-element group 8: 	84 
    -- CP-element group 8: 	208 
    -- CP-element group 8: 	227 
    -- CP-element group 8: 	265 
    -- CP-element group 8: 	246 
    -- CP-element group 8: 	105 
    -- CP-element group 8: 	126 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	276 
    -- CP-element group 9: 	277 
    -- CP-element group 9: 	140 
    -- CP-element group 9: 	181 
    -- CP-element group 9: 	161 
    -- CP-element group 9: 	160 
    -- CP-element group 9: 	182 
    -- CP-element group 9: 	200 
    -- CP-element group 9: 	201 
    -- CP-element group 9: 	293 
    -- CP-element group 9: 	294 
    -- CP-element group 9: 	312 
    -- CP-element group 9: 	313 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	76 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	497 
    -- CP-element group 9: 	498 
    -- CP-element group 9: 	442 
    -- CP-element group 9: 	443 
    -- CP-element group 9: 	219 
    -- CP-element group 9: 	220 
    -- CP-element group 9: 	139 
    -- CP-element group 9: 	388 
    -- CP-element group 9: 	551 
    -- CP-element group 9: 	387 
    -- CP-element group 9: 	238 
    -- CP-element group 9: 	239 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	258 
    -- CP-element group 9: 	332 
    -- CP-element group 9: 	333 
    -- CP-element group 9: 	257 
    -- CP-element group 9: 	97 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	119 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	551 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_42_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(551) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	276 
    -- CP-element group 11: 	181 
    -- CP-element group 11: 	160 
    -- CP-element group 11: 	200 
    -- CP-element group 11: 	293 
    -- CP-element group 11: 	312 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	219 
    -- CP-element group 11: 	139 
    -- CP-element group 11: 	238 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	257 
    -- CP-element group 11: 	97 
    -- CP-element group 11: 	118 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	141 
    -- CP-element group 11: 	162 
    -- CP-element group 11: 	183 
    -- CP-element group 11: 	202 
    -- CP-element group 11: 	295 
    -- CP-element group 11: 	314 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11: 	221 
    -- CP-element group 11: 	240 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	259 
    -- CP-element group 11: 	99 
    -- CP-element group 11: 	120 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= access_T_CP_0_elements(276) & access_T_CP_0_elements(181) & access_T_CP_0_elements(160) & access_T_CP_0_elements(200) & access_T_CP_0_elements(293) & access_T_CP_0_elements(312) & access_T_CP_0_elements(34) & access_T_CP_0_elements(55) & access_T_CP_0_elements(76) & access_T_CP_0_elements(219) & access_T_CP_0_elements(139) & access_T_CP_0_elements(238) & access_T_CP_0_elements(15) & access_T_CP_0_elements(257) & access_T_CP_0_elements(97) & access_T_CP_0_elements(118) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	278 
    -- CP-element group 12: 	142 
    -- CP-element group 12: 	163 
    -- CP-element group 12: 	184 
    -- CP-element group 12: 	296 
    -- CP-element group 12: 	315 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	58 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	203 
    -- CP-element group 12: 	222 
    -- CP-element group 12: 	241 
    -- CP-element group 12: 	260 
    -- CP-element group 12: 	100 
    -- CP-element group 12: 	121 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	552 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	276 
    -- CP-element group 12: 	181 
    -- CP-element group 12: 	160 
    -- CP-element group 12: 	200 
    -- CP-element group 12: 	293 
    -- CP-element group 12: 	312 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	55 
    -- CP-element group 12: 	76 
    -- CP-element group 12: 	219 
    -- CP-element group 12: 	139 
    -- CP-element group 12: 	238 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	257 
    -- CP-element group 12: 	97 
    -- CP-element group 12: 	118 
    -- CP-element group 12:  members (17) 
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= access_T_CP_0_elements(278) & access_T_CP_0_elements(142) & access_T_CP_0_elements(163) & access_T_CP_0_elements(184) & access_T_CP_0_elements(296) & access_T_CP_0_elements(315) & access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(58) & access_T_CP_0_elements(79) & access_T_CP_0_elements(203) & access_T_CP_0_elements(222) & access_T_CP_0_elements(241) & access_T_CP_0_elements(260) & access_T_CP_0_elements(100) & access_T_CP_0_elements(121);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	277 
    -- CP-element group 13: 	140 
    -- CP-element group 13: 	161 
    -- CP-element group 13: 	182 
    -- CP-element group 13: 	201 
    -- CP-element group 13: 	294 
    -- CP-element group 13: 	313 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	77 
    -- CP-element group 13: 	220 
    -- CP-element group 13: 	239 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	258 
    -- CP-element group 13: 	98 
    -- CP-element group 13: 	119 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	143 
    -- CP-element group 13: 	164 
    -- CP-element group 13: 	185 
    -- CP-element group 13: 	297 
    -- CP-element group 13: 	316 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	59 
    -- CP-element group 13: 	80 
    -- CP-element group 13: 	204 
    -- CP-element group 13: 	223 
    -- CP-element group 13: 	242 
    -- CP-element group 13: 	261 
    -- CP-element group 13: 	101 
    -- CP-element group 13: 	122 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= access_T_CP_0_elements(277) & access_T_CP_0_elements(140) & access_T_CP_0_elements(161) & access_T_CP_0_elements(182) & access_T_CP_0_elements(201) & access_T_CP_0_elements(294) & access_T_CP_0_elements(313) & access_T_CP_0_elements(35) & access_T_CP_0_elements(56) & access_T_CP_0_elements(77) & access_T_CP_0_elements(220) & access_T_CP_0_elements(239) & access_T_CP_0_elements(16) & access_T_CP_0_elements(258) & access_T_CP_0_elements(98) & access_T_CP_0_elements(119);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	279 
    -- CP-element group 14: 	144 
    -- CP-element group 14: 	186 
    -- CP-element group 14: 	165 
    -- CP-element group 14: 	298 
    -- CP-element group 14: 	317 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	205 
    -- CP-element group 14: 	224 
    -- CP-element group 14: 	243 
    -- CP-element group 14: 	262 
    -- CP-element group 14: 	102 
    -- CP-element group 14: 	123 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= access_T_CP_0_elements(279) & access_T_CP_0_elements(144) & access_T_CP_0_elements(186) & access_T_CP_0_elements(165) & access_T_CP_0_elements(298) & access_T_CP_0_elements(317) & access_T_CP_0_elements(20) & access_T_CP_0_elements(39) & access_T_CP_0_elements(60) & access_T_CP_0_elements(81) & access_T_CP_0_elements(205) & access_T_CP_0_elements(224) & access_T_CP_0_elements(243) & access_T_CP_0_elements(262) & access_T_CP_0_elements(102) & access_T_CP_0_elements(123);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	367 
    -- CP-element group 16: 	374 
    -- CP-element group 16: 	334 
    -- CP-element group 16: 	360 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(367) & access_T_CP_0_elements(374) & access_T_CP_0_elements(334) & access_T_CP_0_elements(360);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_sample_start__ps
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_update_start__ps
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(13);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	365 
    -- CP-element group 20: 	372 
    -- CP-element group 20: 	14 
    -- CP-element group 20: 	334 
    -- CP-element group 20: 	358 
    -- CP-element group 20:  members (15) 
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_scaled_1
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_resized_1
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_scale_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_scale_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_Sample/req
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_scale_1/scale_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_scale_1/scale_rename_req
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_resize_1/index_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_resize_1/index_resize_req
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_resize_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_resize_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_index_computed_1
      -- 
    req_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => array_obj_ref_138_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_loopback_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_loopback_sample_req_ps
      -- 
    phi_stmt_44_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_44_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_44_req_1); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_entry_trigger
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_entry_sample_req_ps
      -- 
    phi_stmt_44_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_44_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => phi_stmt_44_req_0); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_phi_mux_ack_ps
      -- 
    phi_stmt_44_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_44_ack_0, ack => access_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_update_start_
      -- 
    -- Element group access_T_CP_0_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_update_completed__ps
      -- 
    access_T_CP_0_elements(28) <= access_T_CP_0_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(27), ack => access_T_CP_0_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Sample/req
      -- 
    req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(30), ack => n_address1_210_48_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_update_start_
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Update/req
      -- 
    req_76_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_76_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(31), ack => n_address1_210_48_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Sample/ack
      -- 
    ack_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_210_48_buf_ack_0, ack => access_T_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Update/ack
      -- 
    ack_77_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_210_48_buf_ack_1, ack => access_T_CP_0_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_sample_start_
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	415 
    -- CP-element group 35: 	422 
    -- CP-element group 35: 	429 
    -- CP-element group 35: 	389 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_update_start_
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(415) & access_T_CP_0_elements(422) & access_T_CP_0_elements(429) & access_T_CP_0_elements(389);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_sample_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_update_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(13);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	413 
    -- CP-element group 39: 	420 
    -- CP-element group 39: 	427 
    -- CP-element group 39: 	389 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (15) 
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_resized_1
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_scaled_1
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_computed_1
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_resize_1/$entry
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_resize_1/$exit
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_resize_1/index_resize_req
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_resize_1/index_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_scale_1/$entry
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_scale_1/$exit
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_scale_1/scale_rename_req
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_index_scale_1/scale_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_Sample/req
      -- 
    req_1097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(39), ack => array_obj_ref_311_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_loopback_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_loopback_sample_req_ps
      -- 
    phi_stmt_49_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_49_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_49_req_0); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_entry_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_entry_sample_req_ps
      -- 
    phi_stmt_49_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_49_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_49_req_1); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_phi_mux_ack_ps
      -- 
    phi_stmt_49_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_49_ack_0, ack => access_T_CP_0_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_Sample/req
      -- 
    req_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(45), ack => n_address2_382_51_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_update_start_
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_Update/req
      -- 
    req_112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(46), ack => n_address2_382_51_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_Sample/ack
      -- 
    ack_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_382_51_buf_ack_0, ack => access_T_CP_0_elements(47)); -- 
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_update_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_51_Update/ack
      -- 
    ack_113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_382_51_buf_ack_1, ack => access_T_CP_0_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_Sample/rr
      -- 
    rr_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(51), ack => type_cast_53_inst_req_0); -- 
    access_T_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(49) & access_T_CP_0_elements(53);
      gj_access_T_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_update_start_
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_Update/cr
      -- 
    cr_130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(52), ack => type_cast_53_inst_req_1); -- 
    access_T_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(50) & access_T_CP_0_elements(54);
      gj_access_T_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_Sample/ra
      -- 
    ra_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_53_inst_ack_0, ack => access_T_CP_0_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_53_Update/ca
      -- 
    ca_131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_53_inst_ack_1, ack => access_T_CP_0_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_sample_start_
      -- 
    access_T_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	444 
    -- CP-element group 56: 	470 
    -- CP-element group 56: 	477 
    -- CP-element group 56: 	484 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_update_start_
      -- 
    access_T_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(444) & access_T_CP_0_elements(470) & access_T_CP_0_elements(477) & access_T_CP_0_elements(484);
      gj_access_T_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_sample_start__ps
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_update_start__ps
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(13);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	444 
    -- CP-element group 60: 	475 
    -- CP-element group 60: 	482 
    -- CP-element group 60: 	468 
    -- CP-element group 60: 	14 
    -- CP-element group 60:  members (15) 
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_update_completed__ps
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_resized_1
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_scaled_1
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_computed_1
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_resize_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_resize_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_resize_1/index_resize_req
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_resize_1/index_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_scale_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_scale_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_scale_1/scale_rename_req
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_index_scale_1/scale_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_Sample/req
      -- 
    req_1361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => array_obj_ref_483_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_loopback_trigger
      -- 
    access_T_CP_0_elements(61) <= access_T_CP_0_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_loopback_sample_req_ps
      -- 
    phi_stmt_54_loopback_sample_req_142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_54_loopback_sample_req_142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => phi_stmt_54_req_0); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_entry_trigger
      -- 
    access_T_CP_0_elements(63) <= access_T_CP_0_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_entry_sample_req_ps
      -- 
    phi_stmt_54_entry_sample_req_145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_54_entry_sample_req_145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => phi_stmt_54_req_1); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_phi_mux_ack_ps
      -- 
    phi_stmt_54_phi_mux_ack_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_54_ack_0, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_Sample/req
      -- 
    req_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(66), ack => n_address3_554_56_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_update_start_
      -- CP-element group 67: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_Update/req
      -- 
    req_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(67), ack => n_address3_554_56_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_Sample/ack
      -- 
    ack_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_554_56_buf_ack_0, ack => access_T_CP_0_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_56_Update/ack
      -- 
    ack_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_554_56_buf_ack_1, ack => access_T_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_Sample/rr
      -- 
    rr_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(72), ack => type_cast_58_inst_req_0); -- 
    access_T_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(70) & access_T_CP_0_elements(74);
      gj_access_T_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_update_start_
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_Update/cr
      -- 
    cr_184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(73), ack => type_cast_58_inst_req_1); -- 
    access_T_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(71) & access_T_CP_0_elements(75);
      gj_access_T_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_Sample/ra
      -- 
    ra_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_0, ack => access_T_CP_0_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_58_Update/ca
      -- 
    ca_185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_1, ack => access_T_CP_0_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	9 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	12 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	11 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_sample_start_
      -- 
    access_T_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	499 
    -- CP-element group 77: 	525 
    -- CP-element group 77: 	532 
    -- CP-element group 77: 	539 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_update_start_
      -- 
    access_T_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(499) & access_T_CP_0_elements(525) & access_T_CP_0_elements(532) & access_T_CP_0_elements(539);
      gj_access_T_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	11 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_sample_start__ps
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(11);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	12 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	13 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_update_start__ps
      -- 
    access_T_CP_0_elements(80) <= access_T_CP_0_elements(13);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	499 
    -- CP-element group 81: 	523 
    -- CP-element group 81: 	530 
    -- CP-element group 81: 	537 
    -- CP-element group 81: 	14 
    -- CP-element group 81:  members (15) 
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_update_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_Sample/req
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_scale_1/scale_rename_ack
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_scale_1/scale_rename_req
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_scale_1/$exit
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_scale_1/$entry
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_resize_1/index_resize_ack
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_resize_1/index_resize_req
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_resize_1/$exit
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_resize_1/$entry
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_computed_1
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_scaled_1
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_index_resized_1
      -- 
    req_1625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(81), ack => array_obj_ref_655_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	7 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_loopback_trigger
      -- 
    access_T_CP_0_elements(82) <= access_T_CP_0_elements(7);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_loopback_sample_req_ps
      -- 
    phi_stmt_59_loopback_sample_req_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_59_loopback_sample_req_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => phi_stmt_59_req_1); -- 
    -- Element group access_T_CP_0_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_entry_trigger
      -- 
    access_T_CP_0_elements(84) <= access_T_CP_0_elements(8);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_entry_sample_req_ps
      -- 
    phi_stmt_59_entry_sample_req_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_59_entry_sample_req_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(85), ack => phi_stmt_59_req_0); -- 
    -- Element group access_T_CP_0_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_phi_mux_ack
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_phi_mux_ack_ps
      -- 
    phi_stmt_59_phi_mux_ack_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_59_ack_0, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_Sample/rr
      -- 
    rr_215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(89), ack => type_cast_64_inst_req_0); -- 
    access_T_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(87) & access_T_CP_0_elements(91);
      gj_access_T_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_update_start_
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_Update/cr
      -- 
    cr_220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(90), ack => type_cast_64_inst_req_1); -- 
    access_T_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(88) & access_T_CP_0_elements(92);
      gj_access_T_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_Sample/ra
      -- 
    ra_216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => access_T_CP_0_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_64_Update/ca
      -- 
    ca_221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => access_T_CP_0_elements(92)); -- 
    -- CP-element group 93:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_sample_start__ps
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_Sample/req
      -- 
    req_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(93), ack => n_address4_726_65_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_update_start__ps
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_update_start_
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_Update/req
      -- 
    req_238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(94), ack => n_address4_726_65_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_Sample/ack
      -- 
    ack_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address4_726_65_buf_ack_0, ack => access_T_CP_0_elements(95)); -- 
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_65_Update/ack
      -- 
    ack_239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address4_726_65_buf_ack_1, ack => access_T_CP_0_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	9 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	11 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_sample_start_
      -- 
    access_T_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	367 
    -- CP-element group 98: 	374 
    -- CP-element group 98: 	381 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	13 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_update_start_
      -- 
    access_T_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(367) & access_T_CP_0_elements(374) & access_T_CP_0_elements(381);
      gj_access_T_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	11 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_sample_start__ps
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(11);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	12 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	13 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_update_start__ps
      -- 
    access_T_CP_0_elements(101) <= access_T_CP_0_elements(13);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	365 
    -- CP-element group 102: 	372 
    -- CP-element group 102: 	379 
    -- CP-element group 102: 	14 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	7 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_loopback_trigger
      -- 
    access_T_CP_0_elements(103) <= access_T_CP_0_elements(7);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_loopback_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_loopback_sample_req
      -- 
    phi_stmt_66_loopback_sample_req_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_loopback_sample_req_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(104), ack => phi_stmt_66_req_1); -- 
    -- Element group access_T_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	8 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_entry_trigger
      -- 
    access_T_CP_0_elements(105) <= access_T_CP_0_elements(8);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_entry_sample_req
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_entry_sample_req_ps
      -- 
    phi_stmt_66_entry_sample_req_253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_entry_sample_req_253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(106), ack => phi_stmt_66_req_0); -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_66_phi_mux_ack_ps
      -- 
    phi_stmt_66_phi_mux_ack_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_66_ack_0, ack => access_T_CP_0_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_Sample/rr
      -- 
    rr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(110), ack => type_cast_69_inst_req_0); -- 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(108) & access_T_CP_0_elements(112);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_update_start_
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_Update/cr
      -- 
    cr_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(111), ack => type_cast_69_inst_req_1); -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(109) & access_T_CP_0_elements(113);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_sample_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_Sample/ra
      -- 
    ra_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_0, ack => access_T_CP_0_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_69_Update/ca
      -- 
    ca_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_1, ack => access_T_CP_0_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_Sample/req
      -- 
    req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(114), ack => n_mycounter1_185_70_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_update_start_
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_Update/req
      -- 
    req_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(115), ack => n_mycounter1_185_70_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_sample_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_Sample/ack
      -- 
    ack_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter1_185_70_buf_ack_0, ack => access_T_CP_0_elements(116)); -- 
    -- CP-element group 117:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_update_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_70_Update/ack
      -- 
    ack_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter1_185_70_buf_ack_1, ack => access_T_CP_0_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	12 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	11 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_sample_start_
      -- 
    access_T_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	436 
    -- CP-element group 119: 	422 
    -- CP-element group 119: 	429 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	13 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_update_start_
      -- 
    access_T_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(436) & access_T_CP_0_elements(422) & access_T_CP_0_elements(429);
      gj_access_T_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	11 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_sample_start__ps
      -- 
    access_T_CP_0_elements(120) <= access_T_CP_0_elements(11);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	12 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	13 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_update_start__ps
      -- 
    access_T_CP_0_elements(122) <= access_T_CP_0_elements(13);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	434 
    -- CP-element group 123: 	420 
    -- CP-element group 123: 	427 
    -- CP-element group 123: 	14 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	7 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_loopback_trigger
      -- 
    access_T_CP_0_elements(124) <= access_T_CP_0_elements(7);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_loopback_sample_req
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_loopback_sample_req_ps
      -- 
    phi_stmt_71_loopback_sample_req_304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_loopback_sample_req_304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => phi_stmt_71_req_1); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	8 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_entry_trigger
      -- 
    access_T_CP_0_elements(126) <= access_T_CP_0_elements(8);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_entry_sample_req
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_entry_sample_req_ps
      -- 
    phi_stmt_71_entry_sample_req_307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_entry_sample_req_307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(127), ack => phi_stmt_71_req_0); -- 
    -- Element group access_T_CP_0_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_phi_mux_ack
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_71_phi_mux_ack_ps
      -- 
    phi_stmt_71_phi_mux_ack_310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_71_ack_0, ack => access_T_CP_0_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_Sample/rr
      -- 
    rr_323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(131), ack => type_cast_74_inst_req_0); -- 
    access_T_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(129) & access_T_CP_0_elements(133);
      gj_access_T_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_update_start_
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_Update/cr
      -- 
    cr_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(132), ack => type_cast_74_inst_req_1); -- 
    access_T_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(130) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_Sample/ra
      -- 
    ra_324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_74_inst_ack_0, ack => access_T_CP_0_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_74_Update/ca
      -- 
    ca_329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_74_inst_ack_1, ack => access_T_CP_0_elements(134)); -- 
    -- CP-element group 135:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_sample_start__ps
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_Sample/req
      -- 
    req_341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(135), ack => n_mycounter2_357_75_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_update_start__ps
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_update_start_
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_Update/req
      -- 
    req_346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => n_mycounter2_357_75_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_sample_completed__ps
      -- CP-element group 137: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_Sample/ack
      -- 
    ack_342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter2_357_75_buf_ack_0, ack => access_T_CP_0_elements(137)); -- 
    -- CP-element group 138:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_update_completed__ps
      -- CP-element group 138: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_75_Update/ack
      -- 
    ack_347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter2_357_75_buf_ack_1, ack => access_T_CP_0_elements(138)); -- 
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	9 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	12 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	11 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_sample_start_
      -- 
    access_T_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	9 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	477 
    -- CP-element group 140: 	484 
    -- CP-element group 140: 	491 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	13 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_update_start_
      -- 
    access_T_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(477) & access_T_CP_0_elements(484) & access_T_CP_0_elements(491);
      gj_access_T_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	11 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_sample_start__ps
      -- 
    access_T_CP_0_elements(141) <= access_T_CP_0_elements(11);
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	12 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	13 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_update_start__ps
      -- 
    access_T_CP_0_elements(143) <= access_T_CP_0_elements(13);
    -- CP-element group 144:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	475 
    -- CP-element group 144: 	482 
    -- CP-element group 144: 	489 
    -- CP-element group 144: 	14 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	7 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_loopback_trigger
      -- 
    access_T_CP_0_elements(145) <= access_T_CP_0_elements(7);
    -- CP-element group 146:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_loopback_sample_req
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_loopback_sample_req_ps
      -- 
    phi_stmt_76_loopback_sample_req_358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_loopback_sample_req_358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(146), ack => phi_stmt_76_req_1); -- 
    -- Element group access_T_CP_0_elements(146) is bound as output of CP function.
    -- CP-element group 147:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	8 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_entry_trigger
      -- 
    access_T_CP_0_elements(147) <= access_T_CP_0_elements(8);
    -- CP-element group 148:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_entry_sample_req
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_entry_sample_req_ps
      -- 
    phi_stmt_76_entry_sample_req_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_entry_sample_req_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => phi_stmt_76_req_0); -- 
    -- Element group access_T_CP_0_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_phi_mux_ack
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_76_phi_mux_ack_ps
      -- 
    phi_stmt_76_phi_mux_ack_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_76_ack_0, ack => access_T_CP_0_elements(149)); -- 
    -- CP-element group 150:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (1) 
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_Sample/rr
      -- 
    rr_377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(152), ack => type_cast_79_inst_req_0); -- 
    access_T_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(150) & access_T_CP_0_elements(154);
      gj_access_T_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_update_start_
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_Update/cr
      -- 
    cr_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(153), ack => type_cast_79_inst_req_1); -- 
    access_T_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(151) & access_T_CP_0_elements(155);
      gj_access_T_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_sample_completed__ps
      -- CP-element group 154: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_Sample/ra
      -- 
    ra_378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_79_inst_ack_0, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_update_completed__ps
      -- CP-element group 155: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_79_Update/ca
      -- 
    ca_383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_79_inst_ack_1, ack => access_T_CP_0_elements(155)); -- 
    -- CP-element group 156:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (4) 
      -- CP-element group 156: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_sample_start__ps
      -- CP-element group 156: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_Sample/req
      -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => n_mycounter3_529_80_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(156) is bound as output of CP function.
    -- CP-element group 157:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (4) 
      -- CP-element group 157: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_update_start__ps
      -- CP-element group 157: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_update_start_
      -- CP-element group 157: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_Update/req
      -- 
    req_400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(157), ack => n_mycounter3_529_80_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(157) is bound as output of CP function.
    -- CP-element group 158:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (4) 
      -- CP-element group 158: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_sample_completed__ps
      -- CP-element group 158: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_Sample/ack
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter3_529_80_buf_ack_0, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (4) 
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_update_completed__ps
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_80_Update/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter3_529_80_buf_ack_1, ack => access_T_CP_0_elements(159)); -- 
    -- CP-element group 160:  join  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	9 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	12 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	11 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_sample_start_
      -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	9 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	532 
    -- CP-element group 161: 	539 
    -- CP-element group 161: 	546 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	13 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_update_start_
      -- 
    access_T_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(532) & access_T_CP_0_elements(539) & access_T_CP_0_elements(546);
      gj_access_T_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	11 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_sample_start__ps
      -- 
    access_T_CP_0_elements(162) <= access_T_CP_0_elements(11);
    -- CP-element group 163:  join  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	12 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(163) is bound as output of CP function.
    -- CP-element group 164:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	13 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_update_start__ps
      -- 
    access_T_CP_0_elements(164) <= access_T_CP_0_elements(13);
    -- CP-element group 165:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	530 
    -- CP-element group 165: 	537 
    -- CP-element group 165: 	544 
    -- CP-element group 165: 	14 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(165) is bound as output of CP function.
    -- CP-element group 166:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	7 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_loopback_trigger
      -- 
    access_T_CP_0_elements(166) <= access_T_CP_0_elements(7);
    -- CP-element group 167:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_loopback_sample_req
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_loopback_sample_req_ps
      -- 
    phi_stmt_81_loopback_sample_req_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_81_loopback_sample_req_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => phi_stmt_81_req_1); -- 
    -- Element group access_T_CP_0_elements(167) is bound as output of CP function.
    -- CP-element group 168:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	8 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_entry_trigger
      -- 
    access_T_CP_0_elements(168) <= access_T_CP_0_elements(8);
    -- CP-element group 169:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_entry_sample_req
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_entry_sample_req_ps
      -- 
    phi_stmt_81_entry_sample_req_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_81_entry_sample_req_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(169), ack => phi_stmt_81_req_0); -- 
    -- Element group access_T_CP_0_elements(169) is bound as output of CP function.
    -- CP-element group 170:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (2) 
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_phi_mux_ack
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_81_phi_mux_ack_ps
      -- 
    phi_stmt_81_phi_mux_ack_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_81_ack_0, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(171) is bound as output of CP function.
    -- CP-element group 172:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (1) 
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(172) is bound as output of CP function.
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_Sample/rr
      -- 
    rr_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(173), ack => type_cast_84_inst_req_0); -- 
    access_T_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(171) & access_T_CP_0_elements(175);
      gj_access_T_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_update_start_
      -- CP-element group 174: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_Update/cr
      -- 
    cr_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(174), ack => type_cast_84_inst_req_1); -- 
    access_T_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(172) & access_T_CP_0_elements(176);
      gj_access_T_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (4) 
      -- CP-element group 175: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_sample_completed__ps
      -- CP-element group 175: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_Sample/ra
      -- 
    ra_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_84_inst_ack_0, ack => access_T_CP_0_elements(175)); -- 
    -- CP-element group 176:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (4) 
      -- CP-element group 176: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_update_completed__ps
      -- CP-element group 176: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_84_Update/ca
      -- 
    ca_437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_84_inst_ack_1, ack => access_T_CP_0_elements(176)); -- 
    -- CP-element group 177:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (4) 
      -- CP-element group 177: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_sample_start__ps
      -- CP-element group 177: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_Sample/req
      -- 
    req_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(177), ack => n_mycounter4_701_85_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(177) is bound as output of CP function.
    -- CP-element group 178:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (4) 
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_update_start__ps
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_update_start_
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_Update/req
      -- 
    req_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(178), ack => n_mycounter4_701_85_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(178) is bound as output of CP function.
    -- CP-element group 179:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (4) 
      -- CP-element group 179: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_sample_completed__ps
      -- CP-element group 179: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_Sample/ack
      -- 
    ack_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter4_701_85_buf_ack_0, ack => access_T_CP_0_elements(179)); -- 
    -- CP-element group 180:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (4) 
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_update_completed__ps
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_85_Update/ack
      -- 
    ack_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter4_701_85_buf_ack_1, ack => access_T_CP_0_elements(180)); -- 
    -- CP-element group 181:  join  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	9 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	12 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	11 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_sample_start_
      -- 
    access_T_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	9 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	367 
    -- CP-element group 182: 	374 
    -- CP-element group 182: 	381 
    -- CP-element group 182: 	360 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	13 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_update_start_
      -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(367) & access_T_CP_0_elements(374) & access_T_CP_0_elements(381) & access_T_CP_0_elements(360);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	11 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_sample_start__ps
      -- 
    access_T_CP_0_elements(183) <= access_T_CP_0_elements(11);
    -- CP-element group 184:  join  transition  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	12 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(184) is bound as output of CP function.
    -- CP-element group 185:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	13 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_update_start__ps
      -- 
    access_T_CP_0_elements(185) <= access_T_CP_0_elements(13);
    -- CP-element group 186:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	365 
    -- CP-element group 186: 	372 
    -- CP-element group 186: 	379 
    -- CP-element group 186: 	14 
    -- CP-element group 186: 	358 
    -- CP-element group 186:  members (2) 
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(186) is bound as output of CP function.
    -- CP-element group 187:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	7 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_loopback_trigger
      -- 
    access_T_CP_0_elements(187) <= access_T_CP_0_elements(7);
    -- CP-element group 188:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (2) 
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_loopback_sample_req
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_loopback_sample_req_ps
      -- 
    phi_stmt_86_loopback_sample_req_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_86_loopback_sample_req_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(188), ack => phi_stmt_86_req_0); -- 
    -- Element group access_T_CP_0_elements(188) is bound as output of CP function.
    -- CP-element group 189:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	8 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (1) 
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_entry_trigger
      -- 
    access_T_CP_0_elements(189) <= access_T_CP_0_elements(8);
    -- CP-element group 190:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_entry_sample_req
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_entry_sample_req_ps
      -- 
    phi_stmt_86_entry_sample_req_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_86_entry_sample_req_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => phi_stmt_86_req_1); -- 
    -- Element group access_T_CP_0_elements(190) is bound as output of CP function.
    -- CP-element group 191:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (2) 
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_phi_mux_ack
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_86_phi_mux_ack_ps
      -- 
    phi_stmt_86_phi_mux_ack_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_86_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (4) 
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_sample_start__ps
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_Sample/req
      -- 
    req_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(192), ack => n_row1_193_88_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(192) is bound as output of CP function.
    -- CP-element group 193:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (4) 
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_update_start__ps
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_update_start_
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_Update/req
      -- 
    req_490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => n_row1_193_88_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(193) is bound as output of CP function.
    -- CP-element group 194:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (4) 
      -- CP-element group 194: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_sample_completed__ps
      -- CP-element group 194: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_Sample/ack
      -- 
    ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_193_88_buf_ack_0, ack => access_T_CP_0_elements(194)); -- 
    -- CP-element group 195:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (4) 
      -- CP-element group 195: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_update_completed__ps
      -- CP-element group 195: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_88_Update/ack
      -- 
    ack_491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_193_88_buf_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (4) 
      -- CP-element group 196: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_90_sample_start__ps
      -- CP-element group 196: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_90_sample_completed__ps
      -- CP-element group 196: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_90_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_90_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(196) is bound as output of CP function.
    -- CP-element group 197:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_90_update_start__ps
      -- CP-element group 197: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_90_update_start_
      -- 
    -- Element group access_T_CP_0_elements(197) is bound as output of CP function.
    -- CP-element group 198:  join  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_90_update_completed__ps
      -- 
    access_T_CP_0_elements(198) <= access_T_CP_0_elements(199);
    -- CP-element group 199:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	198 
    -- CP-element group 199:  members (1) 
      -- CP-element group 199: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_90_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(199) is a control-delay.
    cp_element_199_delay: control_delay_element  generic map(name => " 199_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(197), ack => access_T_CP_0_elements(199), clk => clk, reset =>reset);
    -- CP-element group 200:  join  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	9 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	12 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	11 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_sample_start_
      -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  join  transition  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	9 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	436 
    -- CP-element group 201: 	415 
    -- CP-element group 201: 	422 
    -- CP-element group 201: 	429 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	13 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_update_start_
      -- 
    access_T_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(436) & access_T_CP_0_elements(415) & access_T_CP_0_elements(422) & access_T_CP_0_elements(429);
      gj_access_T_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	11 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_sample_start__ps
      -- 
    access_T_CP_0_elements(202) <= access_T_CP_0_elements(11);
    -- CP-element group 203:  join  transition  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	12 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(203) is bound as output of CP function.
    -- CP-element group 204:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	13 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_update_start__ps
      -- 
    access_T_CP_0_elements(204) <= access_T_CP_0_elements(13);
    -- CP-element group 205:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	434 
    -- CP-element group 205: 	413 
    -- CP-element group 205: 	420 
    -- CP-element group 205: 	427 
    -- CP-element group 205: 	14 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(205) is bound as output of CP function.
    -- CP-element group 206:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	7 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_loopback_trigger
      -- 
    access_T_CP_0_elements(206) <= access_T_CP_0_elements(7);
    -- CP-element group 207:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (2) 
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_loopback_sample_req
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_loopback_sample_req_ps
      -- 
    phi_stmt_91_loopback_sample_req_510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_91_loopback_sample_req_510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(207), ack => phi_stmt_91_req_1); -- 
    -- Element group access_T_CP_0_elements(207) is bound as output of CP function.
    -- CP-element group 208:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	8 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (1) 
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_entry_trigger
      -- 
    access_T_CP_0_elements(208) <= access_T_CP_0_elements(8);
    -- CP-element group 209:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (2) 
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_entry_sample_req
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_entry_sample_req_ps
      -- 
    phi_stmt_91_entry_sample_req_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_91_entry_sample_req_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(209), ack => phi_stmt_91_req_0); -- 
    -- Element group access_T_CP_0_elements(209) is bound as output of CP function.
    -- CP-element group 210:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (2) 
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_phi_mux_ack
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_91_phi_mux_ack_ps
      -- 
    phi_stmt_91_phi_mux_ack_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_91_ack_0, ack => access_T_CP_0_elements(210)); -- 
    -- CP-element group 211:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (4) 
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_94_sample_start__ps
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_94_sample_completed__ps
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_94_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_94_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(211) is bound as output of CP function.
    -- CP-element group 212:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (2) 
      -- CP-element group 212: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_94_update_start_
      -- CP-element group 212: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_94_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(212) is bound as output of CP function.
    -- CP-element group 213:  join  transition  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	214 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_94_update_completed__ps
      -- 
    access_T_CP_0_elements(213) <= access_T_CP_0_elements(214);
    -- CP-element group 214:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	213 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_94_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(214) is a control-delay.
    cp_element_214_delay: control_delay_element  generic map(name => " 214_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(212), ack => access_T_CP_0_elements(214), clk => clk, reset =>reset);
    -- CP-element group 215:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (4) 
      -- CP-element group 215: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_sample_start__ps
      -- CP-element group 215: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_Sample/req
      -- 
    req_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(215), ack => n_row2_365_95_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(215) is bound as output of CP function.
    -- CP-element group 216:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (4) 
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_update_start__ps
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_update_start_
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_Update/req
      -- 
    req_542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(216), ack => n_row2_365_95_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(216) is bound as output of CP function.
    -- CP-element group 217:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (4) 
      -- CP-element group 217: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_sample_completed__ps
      -- CP-element group 217: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_Sample/ack
      -- 
    ack_538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_365_95_buf_ack_0, ack => access_T_CP_0_elements(217)); -- 
    -- CP-element group 218:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (4) 
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_update_completed__ps
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_95_Update/ack
      -- 
    ack_543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_365_95_buf_ack_1, ack => access_T_CP_0_elements(218)); -- 
    -- CP-element group 219:  join  transition  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	9 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	12 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	11 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_sample_start_
      -- 
    access_T_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  join  transition  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	9 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	470 
    -- CP-element group 220: 	477 
    -- CP-element group 220: 	484 
    -- CP-element group 220: 	491 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	13 
    -- CP-element group 220:  members (1) 
      -- CP-element group 220: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_update_start_
      -- 
    access_T_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(470) & access_T_CP_0_elements(477) & access_T_CP_0_elements(484) & access_T_CP_0_elements(491);
      gj_access_T_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	11 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (1) 
      -- CP-element group 221: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_sample_start__ps
      -- 
    access_T_CP_0_elements(221) <= access_T_CP_0_elements(11);
    -- CP-element group 222:  join  transition  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	12 
    -- CP-element group 222:  members (1) 
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(222) is bound as output of CP function.
    -- CP-element group 223:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	13 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_update_start__ps
      -- 
    access_T_CP_0_elements(223) <= access_T_CP_0_elements(13);
    -- CP-element group 224:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	475 
    -- CP-element group 224: 	482 
    -- CP-element group 224: 	489 
    -- CP-element group 224: 	468 
    -- CP-element group 224: 	14 
    -- CP-element group 224:  members (2) 
      -- CP-element group 224: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(224) is bound as output of CP function.
    -- CP-element group 225:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	7 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_loopback_trigger
      -- 
    access_T_CP_0_elements(225) <= access_T_CP_0_elements(7);
    -- CP-element group 226:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_loopback_sample_req
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_loopback_sample_req_ps
      -- 
    phi_stmt_96_loopback_sample_req_554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_96_loopback_sample_req_554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(226), ack => phi_stmt_96_req_1); -- 
    -- Element group access_T_CP_0_elements(226) is bound as output of CP function.
    -- CP-element group 227:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	8 
    -- CP-element group 227: successors 
    -- CP-element group 227:  members (1) 
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_entry_trigger
      -- 
    access_T_CP_0_elements(227) <= access_T_CP_0_elements(8);
    -- CP-element group 228:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_entry_sample_req
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_entry_sample_req_ps
      -- 
    phi_stmt_96_entry_sample_req_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_96_entry_sample_req_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(228), ack => phi_stmt_96_req_0); -- 
    -- Element group access_T_CP_0_elements(228) is bound as output of CP function.
    -- CP-element group 229:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (2) 
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_phi_mux_ack
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_96_phi_mux_ack_ps
      -- 
    phi_stmt_96_phi_mux_ack_560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_96_ack_0, ack => access_T_CP_0_elements(229)); -- 
    -- CP-element group 230:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (4) 
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_99_sample_start__ps
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_99_sample_completed__ps
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_99_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_99_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(230) is bound as output of CP function.
    -- CP-element group 231:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	233 
    -- CP-element group 231:  members (2) 
      -- CP-element group 231: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_99_update_start__ps
      -- CP-element group 231: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_99_update_start_
      -- 
    -- Element group access_T_CP_0_elements(231) is bound as output of CP function.
    -- CP-element group 232:  join  transition  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	233 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_99_update_completed__ps
      -- 
    access_T_CP_0_elements(232) <= access_T_CP_0_elements(233);
    -- CP-element group 233:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	232 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_99_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(233) is a control-delay.
    cp_element_233_delay: control_delay_element  generic map(name => " 233_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(231), ack => access_T_CP_0_elements(233), clk => clk, reset =>reset);
    -- CP-element group 234:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (4) 
      -- CP-element group 234: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_sample_start__ps
      -- CP-element group 234: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_Sample/req
      -- 
    req_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(234), ack => n_row3_537_100_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(234) is bound as output of CP function.
    -- CP-element group 235:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (4) 
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_update_start__ps
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_update_start_
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_Update/req
      -- 
    req_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(235), ack => n_row3_537_100_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(235) is bound as output of CP function.
    -- CP-element group 236:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (4) 
      -- CP-element group 236: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_sample_completed__ps
      -- CP-element group 236: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_Sample/ack
      -- 
    ack_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row3_537_100_buf_ack_0, ack => access_T_CP_0_elements(236)); -- 
    -- CP-element group 237:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (4) 
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_update_completed__ps
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_100_Update/ack
      -- 
    ack_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row3_537_100_buf_ack_1, ack => access_T_CP_0_elements(237)); -- 
    -- CP-element group 238:  join  transition  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	9 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	12 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	11 
    -- CP-element group 238:  members (1) 
      -- CP-element group 238: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_sample_start_
      -- 
    access_T_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  join  transition  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	9 
    -- CP-element group 239: marked-predecessors 
    -- CP-element group 239: 	525 
    -- CP-element group 239: 	532 
    -- CP-element group 239: 	539 
    -- CP-element group 239: 	546 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	13 
    -- CP-element group 239:  members (1) 
      -- CP-element group 239: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_update_start_
      -- 
    access_T_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(525) & access_T_CP_0_elements(532) & access_T_CP_0_elements(539) & access_T_CP_0_elements(546);
      gj_access_T_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	11 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (1) 
      -- CP-element group 240: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_sample_start__ps
      -- 
    access_T_CP_0_elements(240) <= access_T_CP_0_elements(11);
    -- CP-element group 241:  join  transition  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	12 
    -- CP-element group 241:  members (1) 
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(241) is bound as output of CP function.
    -- CP-element group 242:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	13 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (1) 
      -- CP-element group 242: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_update_start__ps
      -- 
    access_T_CP_0_elements(242) <= access_T_CP_0_elements(13);
    -- CP-element group 243:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	523 
    -- CP-element group 243: 	530 
    -- CP-element group 243: 	537 
    -- CP-element group 243: 	544 
    -- CP-element group 243: 	14 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(243) is bound as output of CP function.
    -- CP-element group 244:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	7 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (1) 
      -- CP-element group 244: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_loopback_trigger
      -- 
    access_T_CP_0_elements(244) <= access_T_CP_0_elements(7);
    -- CP-element group 245:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: successors 
    -- CP-element group 245:  members (2) 
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_loopback_sample_req
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_loopback_sample_req_ps
      -- 
    phi_stmt_101_loopback_sample_req_598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_101_loopback_sample_req_598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(245), ack => phi_stmt_101_req_1); -- 
    -- Element group access_T_CP_0_elements(245) is bound as output of CP function.
    -- CP-element group 246:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	8 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (1) 
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_entry_trigger
      -- 
    access_T_CP_0_elements(246) <= access_T_CP_0_elements(8);
    -- CP-element group 247:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (2) 
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_entry_sample_req
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_entry_sample_req_ps
      -- 
    phi_stmt_101_entry_sample_req_601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_101_entry_sample_req_601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(247), ack => phi_stmt_101_req_0); -- 
    -- Element group access_T_CP_0_elements(247) is bound as output of CP function.
    -- CP-element group 248:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (2) 
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_phi_mux_ack
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_101_phi_mux_ack_ps
      -- 
    phi_stmt_101_phi_mux_ack_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_101_ack_0, ack => access_T_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (4) 
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_104_sample_start__ps
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_104_sample_completed__ps
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_104_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_104_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(249) is bound as output of CP function.
    -- CP-element group 250:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_104_update_start__ps
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_104_update_start_
      -- 
    -- Element group access_T_CP_0_elements(250) is bound as output of CP function.
    -- CP-element group 251:  join  transition  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	252 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (1) 
      -- CP-element group 251: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_104_update_completed__ps
      -- 
    access_T_CP_0_elements(251) <= access_T_CP_0_elements(252);
    -- CP-element group 252:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	251 
    -- CP-element group 252:  members (1) 
      -- CP-element group 252: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_104_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(252) is a control-delay.
    cp_element_252_delay: control_delay_element  generic map(name => " 252_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(250), ack => access_T_CP_0_elements(252), clk => clk, reset =>reset);
    -- CP-element group 253:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (4) 
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_sample_start__ps
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_Sample/req
      -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(253), ack => n_row4_709_105_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(253) is bound as output of CP function.
    -- CP-element group 254:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (4) 
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_update_start__ps
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_update_start_
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_Update/req
      -- 
    req_630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(254), ack => n_row4_709_105_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(254) is bound as output of CP function.
    -- CP-element group 255:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (4) 
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_sample_completed__ps
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_Sample/ack
      -- 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row4_709_105_buf_ack_0, ack => access_T_CP_0_elements(255)); -- 
    -- CP-element group 256:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (4) 
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_update_completed__ps
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_105_Update/ack
      -- 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row4_709_105_buf_ack_1, ack => access_T_CP_0_elements(256)); -- 
    -- CP-element group 257:  join  transition  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	9 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	12 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	11 
    -- CP-element group 257:  members (1) 
      -- CP-element group 257: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_sample_start_
      -- 
    access_T_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	9 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	367 
    -- CP-element group 258: 	374 
    -- CP-element group 258: 	381 
    -- CP-element group 258: 	360 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	13 
    -- CP-element group 258:  members (1) 
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_update_start_
      -- 
    access_T_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(367) & access_T_CP_0_elements(374) & access_T_CP_0_elements(381) & access_T_CP_0_elements(360);
      gj_access_T_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	11 
    -- CP-element group 259: successors 
    -- CP-element group 259:  members (1) 
      -- CP-element group 259: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_sample_start__ps
      -- 
    access_T_CP_0_elements(259) <= access_T_CP_0_elements(11);
    -- CP-element group 260:  join  transition  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	12 
    -- CP-element group 260:  members (1) 
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(260) is bound as output of CP function.
    -- CP-element group 261:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	13 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (1) 
      -- CP-element group 261: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_update_start__ps
      -- 
    access_T_CP_0_elements(261) <= access_T_CP_0_elements(13);
    -- CP-element group 262:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	365 
    -- CP-element group 262: 	372 
    -- CP-element group 262: 	379 
    -- CP-element group 262: 	14 
    -- CP-element group 262: 	358 
    -- CP-element group 262:  members (2) 
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(262) is bound as output of CP function.
    -- CP-element group 263:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	7 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (1) 
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_loopback_trigger
      -- 
    access_T_CP_0_elements(263) <= access_T_CP_0_elements(7);
    -- CP-element group 264:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (2) 
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_loopback_sample_req
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_loopback_sample_req_ps
      -- 
    phi_stmt_106_loopback_sample_req_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_106_loopback_sample_req_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(264), ack => phi_stmt_106_req_1); -- 
    -- Element group access_T_CP_0_elements(264) is bound as output of CP function.
    -- CP-element group 265:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	8 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (1) 
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_entry_trigger
      -- 
    access_T_CP_0_elements(265) <= access_T_CP_0_elements(8);
    -- CP-element group 266:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_entry_sample_req
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_entry_sample_req_ps
      -- 
    phi_stmt_106_entry_sample_req_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_106_entry_sample_req_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(266), ack => phi_stmt_106_req_0); -- 
    -- Element group access_T_CP_0_elements(266) is bound as output of CP function.
    -- CP-element group 267:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (2) 
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_phi_mux_ack
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_106_phi_mux_ack_ps
      -- 
    phi_stmt_106_phi_mux_ack_648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_106_ack_0, ack => access_T_CP_0_elements(267)); -- 
    -- CP-element group 268:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: successors 
    -- CP-element group 268:  members (4) 
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_sample_start__ps
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_sample_completed__ps
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(268) is bound as output of CP function.
    -- CP-element group 269:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (2) 
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_update_start__ps
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_update_start_
      -- 
    -- Element group access_T_CP_0_elements(269) is bound as output of CP function.
    -- CP-element group 270:  join  transition  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	271 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (1) 
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_update_completed__ps
      -- 
    access_T_CP_0_elements(270) <= access_T_CP_0_elements(271);
    -- CP-element group 271:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	270 
    -- CP-element group 271:  members (1) 
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(271) is a control-delay.
    cp_element_271_delay: control_delay_element  generic map(name => " 271_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(269), ack => access_T_CP_0_elements(271), clk => clk, reset =>reset);
    -- CP-element group 272:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (4) 
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_sample_start__ps
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_Sample/req
      -- 
    req_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(272), ack => n_start1_168_110_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(272) is bound as output of CP function.
    -- CP-element group 273:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (4) 
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_update_start__ps
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_update_start_
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_Update/req
      -- 
    req_674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(273), ack => n_start1_168_110_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(273) is bound as output of CP function.
    -- CP-element group 274:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274:  members (4) 
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_sample_completed__ps
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_Sample/ack
      -- 
    ack_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start1_168_110_buf_ack_0, ack => access_T_CP_0_elements(274)); -- 
    -- CP-element group 275:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (4) 
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_update_completed__ps
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_110_Update/ack
      -- 
    ack_675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start1_168_110_buf_ack_1, ack => access_T_CP_0_elements(275)); -- 
    -- CP-element group 276:  join  transition  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	9 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	12 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	11 
    -- CP-element group 276:  members (1) 
      -- CP-element group 276: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_sample_start_
      -- 
    access_T_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  join  transition  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	9 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	436 
    -- CP-element group 277: 	415 
    -- CP-element group 277: 	422 
    -- CP-element group 277: 	429 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	13 
    -- CP-element group 277:  members (1) 
      -- CP-element group 277: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_update_start_
      -- 
    access_T_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(436) & access_T_CP_0_elements(415) & access_T_CP_0_elements(422) & access_T_CP_0_elements(429);
      gj_access_T_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  join  transition  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	12 
    -- CP-element group 278:  members (1) 
      -- CP-element group 278: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(278) is bound as output of CP function.
    -- CP-element group 279:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	434 
    -- CP-element group 279: 	413 
    -- CP-element group 279: 	420 
    -- CP-element group 279: 	427 
    -- CP-element group 279: 	14 
    -- CP-element group 279:  members (2) 
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(279) is bound as output of CP function.
    -- CP-element group 280:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	7 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_loopback_trigger
      -- 
    access_T_CP_0_elements(280) <= access_T_CP_0_elements(7);
    -- CP-element group 281:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_loopback_sample_req
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_loopback_sample_req_ps
      -- 
    phi_stmt_111_loopback_sample_req_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_111_loopback_sample_req_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(281), ack => phi_stmt_111_req_1); -- 
    -- Element group access_T_CP_0_elements(281) is bound as output of CP function.
    -- CP-element group 282:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	8 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_entry_trigger
      -- 
    access_T_CP_0_elements(282) <= access_T_CP_0_elements(8);
    -- CP-element group 283:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (2) 
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_entry_sample_req
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_entry_sample_req_ps
      -- 
    phi_stmt_111_entry_sample_req_689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_111_entry_sample_req_689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(283), ack => phi_stmt_111_req_0); -- 
    -- Element group access_T_CP_0_elements(283) is bound as output of CP function.
    -- CP-element group 284:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: successors 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_phi_mux_ack
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_phi_mux_ack_ps
      -- 
    phi_stmt_111_phi_mux_ack_692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_111_ack_0, ack => access_T_CP_0_elements(284)); -- 
    -- CP-element group 285:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: successors 
    -- CP-element group 285:  members (4) 
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_114_sample_start__ps
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_114_sample_completed__ps
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_114_sample_start_
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_114_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(285) is bound as output of CP function.
    -- CP-element group 286:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_114_update_start__ps
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_114_update_start_
      -- 
    -- Element group access_T_CP_0_elements(286) is bound as output of CP function.
    -- CP-element group 287:  join  transition  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	288 
    -- CP-element group 287: successors 
    -- CP-element group 287:  members (1) 
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_114_update_completed__ps
      -- 
    access_T_CP_0_elements(287) <= access_T_CP_0_elements(288);
    -- CP-element group 288:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	287 
    -- CP-element group 288:  members (1) 
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_114_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(288) is a control-delay.
    cp_element_288_delay: control_delay_element  generic map(name => " 288_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(286), ack => access_T_CP_0_elements(288), clk => clk, reset =>reset);
    -- CP-element group 289:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (4) 
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_sample_start__ps
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_Sample/req
      -- 
    req_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(289), ack => n_start2_340_115_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(289) is bound as output of CP function.
    -- CP-element group 290:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (4) 
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_update_start__ps
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_update_start_
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_Update/req
      -- 
    req_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(290), ack => n_start2_340_115_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(290) is bound as output of CP function.
    -- CP-element group 291:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (4) 
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_sample_completed__ps
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_Sample/ack
      -- 
    ack_714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start2_340_115_buf_ack_0, ack => access_T_CP_0_elements(291)); -- 
    -- CP-element group 292:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292:  members (4) 
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_update_completed__ps
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_115_Update/ack
      -- 
    ack_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start2_340_115_buf_ack_1, ack => access_T_CP_0_elements(292)); -- 
    -- CP-element group 293:  join  transition  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	9 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	12 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	11 
    -- CP-element group 293:  members (1) 
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_sample_start_
      -- 
    access_T_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	9 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	470 
    -- CP-element group 294: 	477 
    -- CP-element group 294: 	484 
    -- CP-element group 294: 	491 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	13 
    -- CP-element group 294:  members (1) 
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_update_start_
      -- 
    access_T_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(470) & access_T_CP_0_elements(477) & access_T_CP_0_elements(484) & access_T_CP_0_elements(491);
      gj_access_T_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	11 
    -- CP-element group 295: successors 
    -- CP-element group 295:  members (1) 
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_sample_start__ps
      -- 
    access_T_CP_0_elements(295) <= access_T_CP_0_elements(11);
    -- CP-element group 296:  join  transition  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	12 
    -- CP-element group 296:  members (1) 
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(296) is bound as output of CP function.
    -- CP-element group 297:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	13 
    -- CP-element group 297: successors 
    -- CP-element group 297:  members (1) 
      -- CP-element group 297: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_update_start__ps
      -- 
    access_T_CP_0_elements(297) <= access_T_CP_0_elements(13);
    -- CP-element group 298:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	475 
    -- CP-element group 298: 	482 
    -- CP-element group 298: 	489 
    -- CP-element group 298: 	468 
    -- CP-element group 298: 	14 
    -- CP-element group 298:  members (2) 
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_update_completed__ps
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(298) is bound as output of CP function.
    -- CP-element group 299:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	7 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (1) 
      -- CP-element group 299: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_loopback_trigger
      -- 
    access_T_CP_0_elements(299) <= access_T_CP_0_elements(7);
    -- CP-element group 300:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: successors 
    -- CP-element group 300:  members (2) 
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_loopback_sample_req
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_loopback_sample_req_ps
      -- 
    phi_stmt_116_loopback_sample_req_730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_116_loopback_sample_req_730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(300), ack => phi_stmt_116_req_1); -- 
    -- Element group access_T_CP_0_elements(300) is bound as output of CP function.
    -- CP-element group 301:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	8 
    -- CP-element group 301: successors 
    -- CP-element group 301:  members (1) 
      -- CP-element group 301: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_entry_trigger
      -- 
    access_T_CP_0_elements(301) <= access_T_CP_0_elements(8);
    -- CP-element group 302:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: successors 
    -- CP-element group 302:  members (2) 
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_entry_sample_req_ps
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_entry_sample_req
      -- 
    phi_stmt_116_entry_sample_req_733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_116_entry_sample_req_733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(302), ack => phi_stmt_116_req_0); -- 
    -- Element group access_T_CP_0_elements(302) is bound as output of CP function.
    -- CP-element group 303:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: successors 
    -- CP-element group 303:  members (2) 
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_phi_mux_ack_ps
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_phi_mux_ack
      -- 
    phi_stmt_116_phi_mux_ack_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_116_ack_0, ack => access_T_CP_0_elements(303)); -- 
    -- CP-element group 304:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (4) 
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_sample_completed_
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_sample_completed__ps
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(304) is bound as output of CP function.
    -- CP-element group 305:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_update_start__ps
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_update_start_
      -- 
    -- Element group access_T_CP_0_elements(305) is bound as output of CP function.
    -- CP-element group 306:  join  transition  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	307 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (1) 
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_update_completed__ps
      -- 
    access_T_CP_0_elements(306) <= access_T_CP_0_elements(307);
    -- CP-element group 307:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	306 
    -- CP-element group 307:  members (1) 
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(307) is a control-delay.
    cp_element_307_delay: control_delay_element  generic map(name => " 307_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(305), ack => access_T_CP_0_elements(307), clk => clk, reset =>reset);
    -- CP-element group 308:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	310 
    -- CP-element group 308:  members (4) 
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_sample_start__ps
      -- 
    req_757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(308), ack => n_start3_512_120_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(308) is bound as output of CP function.
    -- CP-element group 309:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (4) 
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_update_start_
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_update_start__ps
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_Update/req
      -- 
    req_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(309), ack => n_start3_512_120_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(309) is bound as output of CP function.
    -- CP-element group 310:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	308 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (4) 
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_Sample/ack
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_sample_completed__ps
      -- 
    ack_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start3_512_120_buf_ack_0, ack => access_T_CP_0_elements(310)); -- 
    -- CP-element group 311:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311:  members (4) 
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_update_completed__ps
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_120_Update/ack
      -- 
    ack_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start3_512_120_buf_ack_1, ack => access_T_CP_0_elements(311)); -- 
    -- CP-element group 312:  join  transition  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	9 
    -- CP-element group 312: marked-predecessors 
    -- CP-element group 312: 	12 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	11 
    -- CP-element group 312:  members (1) 
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_sample_start_
      -- 
    access_T_cp_element_group_312: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_312"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_312 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(312), clk => clk, reset => reset); --
    end block;
    -- CP-element group 313:  join  transition  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	9 
    -- CP-element group 313: marked-predecessors 
    -- CP-element group 313: 	525 
    -- CP-element group 313: 	532 
    -- CP-element group 313: 	539 
    -- CP-element group 313: 	546 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	13 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_update_start_
      -- 
    access_T_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(525) & access_T_CP_0_elements(532) & access_T_CP_0_elements(539) & access_T_CP_0_elements(546);
      gj_access_T_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	11 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (1) 
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_sample_start__ps
      -- 
    access_T_CP_0_elements(314) <= access_T_CP_0_elements(11);
    -- CP-element group 315:  join  transition  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	12 
    -- CP-element group 315:  members (1) 
      -- CP-element group 315: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(315) is bound as output of CP function.
    -- CP-element group 316:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	13 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (1) 
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_update_start__ps
      -- 
    access_T_CP_0_elements(316) <= access_T_CP_0_elements(13);
    -- CP-element group 317:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	523 
    -- CP-element group 317: 	530 
    -- CP-element group 317: 	537 
    -- CP-element group 317: 	544 
    -- CP-element group 317: 	14 
    -- CP-element group 317:  members (2) 
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_update_completed_
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(317) is bound as output of CP function.
    -- CP-element group 318:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	7 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (1) 
      -- CP-element group 318: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_loopback_trigger
      -- 
    access_T_CP_0_elements(318) <= access_T_CP_0_elements(7);
    -- CP-element group 319:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: successors 
    -- CP-element group 319:  members (2) 
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_loopback_sample_req
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_loopback_sample_req_ps
      -- 
    phi_stmt_121_loopback_sample_req_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_121_loopback_sample_req_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(319), ack => phi_stmt_121_req_1); -- 
    -- Element group access_T_CP_0_elements(319) is bound as output of CP function.
    -- CP-element group 320:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	8 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (1) 
      -- CP-element group 320: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_entry_trigger
      -- 
    access_T_CP_0_elements(320) <= access_T_CP_0_elements(8);
    -- CP-element group 321:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: successors 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_entry_sample_req_ps
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_entry_sample_req
      -- 
    phi_stmt_121_entry_sample_req_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_121_entry_sample_req_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(321), ack => phi_stmt_121_req_0); -- 
    -- Element group access_T_CP_0_elements(321) is bound as output of CP function.
    -- CP-element group 322:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (2) 
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_phi_mux_ack_ps
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_phi_mux_ack
      -- 
    phi_stmt_121_phi_mux_ack_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_121_ack_0, ack => access_T_CP_0_elements(322)); -- 
    -- CP-element group 323:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: successors 
    -- CP-element group 323:  members (4) 
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_124_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_124_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_124_sample_completed__ps
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_124_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(323) is bound as output of CP function.
    -- CP-element group 324:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (2) 
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_124_update_start_
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_124_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(324) is bound as output of CP function.
    -- CP-element group 325:  join  transition  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	326 
    -- CP-element group 325: successors 
    -- CP-element group 325:  members (1) 
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_124_update_completed__ps
      -- 
    access_T_CP_0_elements(325) <= access_T_CP_0_elements(326);
    -- CP-element group 326:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	325 
    -- CP-element group 326:  members (1) 
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_124_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(326) is a control-delay.
    cp_element_326_delay: control_delay_element  generic map(name => " 326_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(324), ack => access_T_CP_0_elements(326), clk => clk, reset =>reset);
    -- CP-element group 327:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (4) 
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_Sample/req
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_Sample/$entry
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_sample_start_
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_sample_start__ps
      -- 
    req_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(327), ack => n_start4_684_125_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(327) is bound as output of CP function.
    -- CP-element group 328:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	330 
    -- CP-element group 328:  members (4) 
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_Update/req
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_update_start_
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_update_start__ps
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_Update/$entry
      -- 
    req_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(328), ack => n_start4_684_125_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(328) is bound as output of CP function.
    -- CP-element group 329:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: successors 
    -- CP-element group 329:  members (4) 
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_sample_completed__ps
      -- 
    ack_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start4_684_125_buf_ack_0, ack => access_T_CP_0_elements(329)); -- 
    -- CP-element group 330:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	328 
    -- CP-element group 330: successors 
    -- CP-element group 330:  members (4) 
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_Update/ack
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_update_completed__ps
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_125_Update/$exit
      -- 
    ack_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start4_684_125_buf_ack_1, ack => access_T_CP_0_elements(330)); -- 
    -- CP-element group 331:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	335 
    -- CP-element group 331: marked-predecessors 
    -- CP-element group 331: 	336 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	336 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_request/req
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_request/$entry
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_sample_start_
      -- 
    req_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(331), ack => addr_of_139_final_reg_req_0); -- 
    access_T_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(335) & access_T_CP_0_elements(336);
      gj_access_T_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	9 
    -- CP-element group 332: marked-predecessors 
    -- CP-element group 332: 	340 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	337 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_complete/req
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_complete/$entry
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_update_start_
      -- 
    req_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(332), ack => addr_of_139_final_reg_req_1); -- 
    access_T_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(340);
      gj_access_T_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	9 
    -- CP-element group 333: marked-predecessors 
    -- CP-element group 333: 	336 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_Update/req
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_update_start
      -- 
    req_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(333), ack => array_obj_ref_138_index_offset_req_1); -- 
    access_T_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(336);
      gj_access_T_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	20 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	552 
    -- CP-element group 334: marked-successors 
    -- CP-element group 334: 	16 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_Sample/ack
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_sample_complete
      -- 
    ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_138_index_offset_ack_0, ack => access_T_CP_0_elements(334)); -- 
    -- CP-element group 335:  transition  input  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	331 
    -- CP-element group 335:  members (8) 
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_offset_calculated
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_root_address_calculated
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_base_plus_offset/sum_rename_ack
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_base_plus_offset/sum_rename_req
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_base_plus_offset/$exit
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_base_plus_offset/$entry
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_Update/ack
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_138_final_index_sum_regn_Update/$exit
      -- 
    ack_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_138_index_offset_ack_1, ack => access_T_CP_0_elements(335)); -- 
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	331 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	331 
    -- CP-element group 336: 	333 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_request/ack
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_request/$exit
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_sample_completed_
      -- 
    ack_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_139_final_reg_ack_0, ack => access_T_CP_0_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	332 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (19) 
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_word_addrgen/root_register_ack
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_word_addrgen/root_register_req
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_word_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_word_addrgen/$exit
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_word_addrgen/$entry
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_complete/ack
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_complete/$exit
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_139_update_completed_
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_plus_offset/sum_rename_ack
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_plus_offset/sum_rename_req
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_plus_offset/$exit
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_plus_offset/$entry
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_addr_resize/base_resize_ack
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_addr_resize/base_resize_req
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_addr_resize/$exit
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_addr_resize/$entry
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_base_address_resized
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_root_address_calculated
      -- 
    ack_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_139_final_reg_ack_1, ack => access_T_CP_0_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (5) 
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Sample/word_access_start/word_0/rr
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Sample/word_access_start/word_0/$entry
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Sample/word_access_start/$entry
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Sample/$entry
      -- 
    rr_887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(338), ack => ptr_deref_143_load_0_req_0); -- 
    access_T_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(337) & access_T_CP_0_elements(340);
      gj_access_T_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	344 
    -- CP-element group 339: 	348 
    -- CP-element group 339: 	352 
    -- CP-element group 339: 	356 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (5) 
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_update_start_
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/word_access_complete/word_0/cr
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/word_access_complete/word_0/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/word_access_complete/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/$entry
      -- 
    cr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(339), ack => ptr_deref_143_load_0_req_1); -- 
    access_T_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(344) & access_T_CP_0_elements(348) & access_T_CP_0_elements(352) & access_T_CP_0_elements(356);
      gj_access_T_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	332 
    -- CP-element group 340: 	338 
    -- CP-element group 340:  members (5) 
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Sample/word_access_start/word_0/ra
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Sample/word_access_start/word_0/$exit
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Sample/word_access_start/$exit
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Sample/$exit
      -- 
    ra_888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_143_load_0_ack_0, ack => access_T_CP_0_elements(340)); -- 
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341: 	346 
    -- CP-element group 341: 	350 
    -- CP-element group 341: 	354 
    -- CP-element group 341:  members (9) 
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/ptr_deref_143_Merge/merge_ack
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/ptr_deref_143_Merge/merge_req
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/ptr_deref_143_Merge/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/ptr_deref_143_Merge/$entry
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/word_access_complete/word_0/ca
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/word_access_complete/word_0/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/word_access_complete/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_143_update_completed_
      -- 
    ca_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_143_load_0_ack_1, ack => access_T_CP_0_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_Sample/rr
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_sample_start_
      -- 
    rr_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(342), ack => slice_147_inst_req_0); -- 
    access_T_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(341) & access_T_CP_0_elements(344);
      gj_access_T_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	363 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_update_start_
      -- 
    cr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(343), ack => slice_147_inst_req_1); -- 
    access_T_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(363);
      gj_access_T_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	339 
    -- CP-element group 344: 	342 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_Sample/ra
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_sample_completed_
      -- 
    ra_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_147_inst_ack_0, ack => access_T_CP_0_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	362 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_Update/ca
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_147_update_completed_
      -- 
    ca_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_147_inst_ack_1, ack => access_T_CP_0_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	341 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_Sample/rr
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_Sample/$entry
      -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(346), ack => slice_151_inst_req_0); -- 
    access_T_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(341) & access_T_CP_0_elements(348);
      gj_access_T_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	370 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	349 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_Update/cr
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_update_start_
      -- 
    cr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(347), ack => slice_151_inst_req_1); -- 
    access_T_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(370);
      gj_access_T_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348: marked-successors 
    -- CP-element group 348: 	339 
    -- CP-element group 348: 	346 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_Sample/ra
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_Sample/$exit
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_151_inst_ack_0, ack => access_T_CP_0_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	347 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	369 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_Update/ca
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_Update/$exit
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_151_update_completed_
      -- 
    ca_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_151_inst_ack_1, ack => access_T_CP_0_elements(349)); -- 
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	341 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	352 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_Sample/rr
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_sample_start_
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_Sample/$entry
      -- 
    rr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(350), ack => slice_155_inst_req_0); -- 
    access_T_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(341) & access_T_CP_0_elements(352);
      gj_access_T_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: marked-predecessors 
    -- CP-element group 351: 	377 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_Update/cr
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_Update/$entry
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_update_start_
      -- 
    cr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(351), ack => slice_155_inst_req_1); -- 
    access_T_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(377);
      gj_access_T_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	339 
    -- CP-element group 352: 	350 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_Sample/ra
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_sample_completed_
      -- 
    ra_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_155_inst_ack_0, ack => access_T_CP_0_elements(352)); -- 
    -- CP-element group 353:  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	376 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_Update/ca
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_155_update_completed_
      -- 
    ca_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_155_inst_ack_1, ack => access_T_CP_0_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	341 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_Sample/rr
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_Sample/$entry
      -- 
    rr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(354), ack => slice_159_inst_req_0); -- 
    access_T_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(341) & access_T_CP_0_elements(356);
      gj_access_T_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: marked-predecessors 
    -- CP-element group 355: 	384 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_Update/cr
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_update_start_
      -- 
    cr_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(355), ack => slice_159_inst_req_1); -- 
    access_T_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(384);
      gj_access_T_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	339 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_Sample/ra
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_Sample/$exit
      -- 
    ra_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_159_inst_ack_0, ack => access_T_CP_0_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	383 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_Update/ca
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_159_update_completed_
      -- 
    ca_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_159_inst_ack_1, ack => access_T_CP_0_elements(357)); -- 
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	186 
    -- CP-element group 358: 	20 
    -- CP-element group 358: 	262 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_Sample/req
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_Sample/$entry
      -- 
    req_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(358), ack => W_send1_1_272_delayed_14_0_272_inst_req_0); -- 
    access_T_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(186) & access_T_CP_0_elements(20) & access_T_CP_0_elements(262) & access_T_CP_0_elements(360);
      gj_access_T_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: marked-predecessors 
    -- CP-element group 359: 	363 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_Update/req
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_update_start_
      -- 
    req_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(359), ack => W_send1_1_272_delayed_14_0_272_inst_req_1); -- 
    access_T_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(363);
      gj_access_T_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	182 
    -- CP-element group 360: 	16 
    -- CP-element group 360: 	258 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_Sample/ack
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_sample_completed_
      -- 
    ack_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send1_1_272_delayed_14_0_272_inst_ack_0, ack => access_T_CP_0_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_274_Update/ack
      -- 
    ack_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send1_1_272_delayed_14_0_272_inst_ack_1, ack => access_T_CP_0_elements(361)); -- 
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	345 
    -- CP-element group 362: 	361 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	385 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_Sample/req
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_sample_start_
      -- 
    req_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(362), ack => WPIPE_input_pipe1_276_inst_req_0); -- 
    access_T_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(345) & access_T_CP_0_elements(361) & access_T_CP_0_elements(385);
      gj_access_T_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363: marked-successors 
    -- CP-element group 363: 	343 
    -- CP-element group 363: 	359 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_Update/req
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_update_start_
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_sample_completed_
      -- 
    ack_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_276_inst_ack_0, ack => access_T_CP_0_elements(363)); -- 
    req_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(363), ack => WPIPE_input_pipe1_276_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	369 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_Update/ack
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_276_update_completed_
      -- 
    ack_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_276_inst_ack_1, ack => access_T_CP_0_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	186 
    -- CP-element group 365: 	20 
    -- CP-element group 365: 	262 
    -- CP-element group 365: 	102 
    -- CP-element group 365: marked-predecessors 
    -- CP-element group 365: 	367 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	367 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_Sample/req
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_Sample/$entry
      -- 
    req_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(365), ack => W_send2_1_276_delayed_14_0_279_inst_req_0); -- 
    access_T_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(186) & access_T_CP_0_elements(20) & access_T_CP_0_elements(262) & access_T_CP_0_elements(102) & access_T_CP_0_elements(367);
      gj_access_T_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	370 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_update_start_
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_Update/req
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_Update/$entry
      -- 
    req_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(366), ack => W_send2_1_276_delayed_14_0_279_inst_req_1); -- 
    access_T_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(370);
      gj_access_T_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	365 
    -- CP-element group 367: successors 
    -- CP-element group 367: marked-successors 
    -- CP-element group 367: 	182 
    -- CP-element group 367: 	365 
    -- CP-element group 367: 	16 
    -- CP-element group 367: 	258 
    -- CP-element group 367: 	98 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_Sample/ack
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_Sample/$exit
      -- 
    ack_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send2_1_276_delayed_14_0_279_inst_ack_0, ack => access_T_CP_0_elements(367)); -- 
    -- CP-element group 368:  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_Update/ack
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_281_update_completed_
      -- 
    ack_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send2_1_276_delayed_14_0_279_inst_ack_1, ack => access_T_CP_0_elements(368)); -- 
    -- CP-element group 369:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: 	349 
    -- CP-element group 369: 	364 
    -- CP-element group 369: marked-predecessors 
    -- CP-element group 369: 	371 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_Sample/req
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_sample_start_
      -- 
    req_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(369), ack => WPIPE_input_pipe1_283_inst_req_0); -- 
    access_T_cp_element_group_369: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_369"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(368) & access_T_CP_0_elements(349) & access_T_CP_0_elements(364) & access_T_CP_0_elements(371);
      gj_access_T_cp_element_group_369 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(369), clk => clk, reset => reset); --
    end block;
    -- CP-element group 370:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	366 
    -- CP-element group 370: 	347 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_update_start_
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_Update/req
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_Sample/ack
      -- 
    ack_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_283_inst_ack_0, ack => access_T_CP_0_elements(370)); -- 
    req_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(370), ack => WPIPE_input_pipe1_283_inst_req_1); -- 
    -- CP-element group 371:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	376 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	369 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_Update/ack
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_283_Update/$exit
      -- 
    ack_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_283_inst_ack_1, ack => access_T_CP_0_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	186 
    -- CP-element group 372: 	20 
    -- CP-element group 372: 	262 
    -- CP-element group 372: 	102 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_Sample/req
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_Sample/$entry
      -- 
    req_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(372), ack => W_send3_1_280_delayed_14_0_286_inst_req_0); -- 
    access_T_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(186) & access_T_CP_0_elements(20) & access_T_CP_0_elements(262) & access_T_CP_0_elements(102) & access_T_CP_0_elements(374);
      gj_access_T_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: marked-predecessors 
    -- CP-element group 373: 	377 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_Update/req
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_update_start_
      -- 
    req_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(373), ack => W_send3_1_280_delayed_14_0_286_inst_req_1); -- 
    access_T_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(377);
      gj_access_T_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	182 
    -- CP-element group 374: 	372 
    -- CP-element group 374: 	16 
    -- CP-element group 374: 	258 
    -- CP-element group 374: 	98 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_Sample/ack
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_Sample/$exit
      -- 
    ack_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send3_1_280_delayed_14_0_286_inst_ack_0, ack => access_T_CP_0_elements(374)); -- 
    -- CP-element group 375:  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_Update/ack
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_288_update_completed_
      -- 
    ack_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send3_1_280_delayed_14_0_286_inst_ack_1, ack => access_T_CP_0_elements(375)); -- 
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	371 
    -- CP-element group 376: 	375 
    -- CP-element group 376: 	353 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_Sample/req
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_Sample/$entry
      -- 
    req_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(376), ack => WPIPE_input_pipe1_290_inst_req_0); -- 
    access_T_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(371) & access_T_CP_0_elements(375) & access_T_CP_0_elements(353) & access_T_CP_0_elements(378);
      gj_access_T_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377: marked-successors 
    -- CP-element group 377: 	373 
    -- CP-element group 377: 	351 
    -- CP-element group 377:  members (6) 
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_Update/$entry
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_update_start_
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_Sample/ack
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_sample_completed_
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_Update/req
      -- 
    ack_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_290_inst_ack_0, ack => access_T_CP_0_elements(377)); -- 
    req_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(377), ack => WPIPE_input_pipe1_290_inst_req_1); -- 
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	383 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_Update/ack
      -- CP-element group 378: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_290_update_completed_
      -- 
    ack_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_290_inst_ack_1, ack => access_T_CP_0_elements(378)); -- 
    -- CP-element group 379:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	186 
    -- CP-element group 379: 	262 
    -- CP-element group 379: 	102 
    -- CP-element group 379: marked-predecessors 
    -- CP-element group 379: 	381 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_Sample/req
      -- 
    req_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(379), ack => W_send4_1_284_delayed_14_0_293_inst_req_0); -- 
    access_T_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(186) & access_T_CP_0_elements(262) & access_T_CP_0_elements(102) & access_T_CP_0_elements(381);
      gj_access_T_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	384 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_update_start_
      -- CP-element group 380: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_Update/req
      -- 
    req_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(380), ack => W_send4_1_284_delayed_14_0_293_inst_req_1); -- 
    access_T_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(384);
      gj_access_T_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: successors 
    -- CP-element group 381: marked-successors 
    -- CP-element group 381: 	182 
    -- CP-element group 381: 	379 
    -- CP-element group 381: 	258 
    -- CP-element group 381: 	98 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_Sample/ack
      -- CP-element group 381: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_sample_completed_
      -- 
    ack_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send4_1_284_delayed_14_0_293_inst_ack_0, ack => access_T_CP_0_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_295_Update/ack
      -- 
    ack_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send4_1_284_delayed_14_0_293_inst_ack_1, ack => access_T_CP_0_elements(382)); -- 
    -- CP-element group 383:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	378 
    -- CP-element group 383: 	382 
    -- CP-element group 383: 	357 
    -- CP-element group 383: marked-predecessors 
    -- CP-element group 383: 	385 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_Sample/req
      -- 
    req_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(383), ack => WPIPE_input_pipe1_297_inst_req_0); -- 
    access_T_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(378) & access_T_CP_0_elements(382) & access_T_CP_0_elements(357) & access_T_CP_0_elements(385);
      gj_access_T_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384: marked-successors 
    -- CP-element group 384: 	380 
    -- CP-element group 384: 	355 
    -- CP-element group 384:  members (6) 
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_update_start_
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_Sample/ack
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_Update/req
      -- 
    ack_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_297_inst_ack_0, ack => access_T_CP_0_elements(384)); -- 
    req_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(384), ack => WPIPE_input_pipe1_297_inst_req_1); -- 
    -- CP-element group 385:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	552 
    -- CP-element group 385: marked-successors 
    -- CP-element group 385: 	383 
    -- CP-element group 385: 	362 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_297_Update/ack
      -- 
    ack_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_297_inst_ack_1, ack => access_T_CP_0_elements(385)); -- 
    -- CP-element group 386:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	390 
    -- CP-element group 386: marked-predecessors 
    -- CP-element group 386: 	391 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	391 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_sample_start_
      -- CP-element group 386: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_request/$entry
      -- CP-element group 386: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_request/req
      -- 
    req_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(386), ack => addr_of_312_final_reg_req_0); -- 
    access_T_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(390) & access_T_CP_0_elements(391);
      gj_access_T_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	9 
    -- CP-element group 387: marked-predecessors 
    -- CP-element group 387: 	395 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	392 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_update_start_
      -- CP-element group 387: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_complete/$entry
      -- CP-element group 387: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_complete/req
      -- 
    req_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(387), ack => addr_of_312_final_reg_req_1); -- 
    access_T_cp_element_group_387: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_387"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(395);
      gj_access_T_cp_element_group_387 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(387), clk => clk, reset => reset); --
    end block;
    -- CP-element group 388:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	9 
    -- CP-element group 388: marked-predecessors 
    -- CP-element group 388: 	391 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	390 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_update_start
      -- CP-element group 388: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_Update/$entry
      -- CP-element group 388: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_Update/req
      -- 
    req_1102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(388), ack => array_obj_ref_311_index_offset_req_1); -- 
    access_T_cp_element_group_388: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_388"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(391);
      gj_access_T_cp_element_group_388 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 389:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	39 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	552 
    -- CP-element group 389: marked-successors 
    -- CP-element group 389: 	35 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_sample_complete
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_Sample/ack
      -- 
    ack_1098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_311_index_offset_ack_0, ack => access_T_CP_0_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	388 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	386 
    -- CP-element group 390:  members (8) 
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_root_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_offset_calculated
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_final_index_sum_regn_Update/ack
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_base_plus_offset/$entry
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_base_plus_offset/$exit
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_base_plus_offset/sum_rename_req
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_311_base_plus_offset/sum_rename_ack
      -- 
    ack_1103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_311_index_offset_ack_1, ack => access_T_CP_0_elements(390)); -- 
    -- CP-element group 391:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	386 
    -- CP-element group 391: successors 
    -- CP-element group 391: marked-successors 
    -- CP-element group 391: 	388 
    -- CP-element group 391: 	386 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_sample_completed_
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_request/$exit
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_request/ack
      -- 
    ack_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_312_final_reg_ack_0, ack => access_T_CP_0_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	387 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (19) 
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_update_completed_
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_complete/$exit
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_312_complete/ack
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_address_calculated
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_word_address_calculated
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_root_address_calculated
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_address_resized
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_addr_resize/$entry
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_addr_resize/$exit
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_addr_resize/base_resize_req
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_addr_resize/base_resize_ack
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_plus_offset/$entry
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_plus_offset/$exit
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_plus_offset/sum_rename_req
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_base_plus_offset/sum_rename_ack
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_word_addrgen/$entry
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_word_addrgen/$exit
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_word_addrgen/root_register_req
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_word_addrgen/root_register_ack
      -- 
    ack_1118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_312_final_reg_ack_1, ack => access_T_CP_0_elements(392)); -- 
    -- CP-element group 393:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: marked-predecessors 
    -- CP-element group 393: 	395 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	395 
    -- CP-element group 393:  members (5) 
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Sample/word_access_start/$entry
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Sample/word_access_start/word_0/$entry
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Sample/word_access_start/word_0/rr
      -- 
    rr_1151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(393), ack => ptr_deref_316_load_0_req_0); -- 
    access_T_cp_element_group_393: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_393"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(392) & access_T_CP_0_elements(395);
      gj_access_T_cp_element_group_393 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(393), clk => clk, reset => reset); --
    end block;
    -- CP-element group 394:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: marked-predecessors 
    -- CP-element group 394: 	403 
    -- CP-element group 394: 	407 
    -- CP-element group 394: 	411 
    -- CP-element group 394: 	399 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	396 
    -- CP-element group 394:  members (5) 
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_update_start_
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/word_access_complete/$entry
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/word_access_complete/word_0/$entry
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/word_access_complete/word_0/cr
      -- 
    cr_1162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(394), ack => ptr_deref_316_load_0_req_1); -- 
    access_T_cp_element_group_394: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_394"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(403) & access_T_CP_0_elements(407) & access_T_CP_0_elements(411) & access_T_CP_0_elements(399);
      gj_access_T_cp_element_group_394 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(394), clk => clk, reset => reset); --
    end block;
    -- CP-element group 395:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	393 
    -- CP-element group 395: successors 
    -- CP-element group 395: marked-successors 
    -- CP-element group 395: 	393 
    -- CP-element group 395: 	387 
    -- CP-element group 395:  members (5) 
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_sample_completed_
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Sample/word_access_start/$exit
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Sample/word_access_start/word_0/$exit
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Sample/word_access_start/word_0/ra
      -- 
    ra_1152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_316_load_0_ack_0, ack => access_T_CP_0_elements(395)); -- 
    -- CP-element group 396:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	394 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	405 
    -- CP-element group 396: 	409 
    -- CP-element group 396: 	397 
    -- CP-element group 396: 	401 
    -- CP-element group 396:  members (9) 
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_update_completed_
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/word_access_complete/$exit
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/word_access_complete/word_0/$exit
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/word_access_complete/word_0/ca
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/ptr_deref_316_Merge/$entry
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/ptr_deref_316_Merge/$exit
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/ptr_deref_316_Merge/merge_req
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_316_Update/ptr_deref_316_Merge/merge_ack
      -- 
    ca_1163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_316_load_0_ack_1, ack => access_T_CP_0_elements(396)); -- 
    -- CP-element group 397:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: marked-predecessors 
    -- CP-element group 397: 	399 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	399 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_Sample/rr
      -- 
    rr_1176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(397), ack => slice_320_inst_req_0); -- 
    access_T_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(396) & access_T_CP_0_elements(399);
      gj_access_T_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: marked-predecessors 
    -- CP-element group 398: 	418 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	400 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_update_start_
      -- CP-element group 398: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_Update/cr
      -- 
    cr_1181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(398), ack => slice_320_inst_req_1); -- 
    access_T_cp_element_group_398: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_398"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(418);
      gj_access_T_cp_element_group_398 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(398), clk => clk, reset => reset); --
    end block;
    -- CP-element group 399:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	397 
    -- CP-element group 399: successors 
    -- CP-element group 399: marked-successors 
    -- CP-element group 399: 	394 
    -- CP-element group 399: 	397 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_Sample/$exit
      -- CP-element group 399: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_Sample/ra
      -- 
    ra_1177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_320_inst_ack_0, ack => access_T_CP_0_elements(399)); -- 
    -- CP-element group 400:  transition  input  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	398 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	417 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_update_completed_
      -- CP-element group 400: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_320_Update/ca
      -- 
    ca_1182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_320_inst_ack_1, ack => access_T_CP_0_elements(400)); -- 
    -- CP-element group 401:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	396 
    -- CP-element group 401: marked-predecessors 
    -- CP-element group 401: 	403 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	403 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_Sample/rr
      -- 
    rr_1190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(401), ack => slice_324_inst_req_0); -- 
    access_T_cp_element_group_401: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_401"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(396) & access_T_CP_0_elements(403);
      gj_access_T_cp_element_group_401 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(401), clk => clk, reset => reset); --
    end block;
    -- CP-element group 402:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: marked-predecessors 
    -- CP-element group 402: 	425 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_update_start_
      -- CP-element group 402: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_Update/cr
      -- 
    cr_1195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(402), ack => slice_324_inst_req_1); -- 
    access_T_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(425);
      gj_access_T_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	401 
    -- CP-element group 403: successors 
    -- CP-element group 403: marked-successors 
    -- CP-element group 403: 	394 
    -- CP-element group 403: 	401 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_sample_completed_
      -- CP-element group 403: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_Sample/ra
      -- 
    ra_1191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_324_inst_ack_0, ack => access_T_CP_0_elements(403)); -- 
    -- CP-element group 404:  transition  input  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	424 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_update_completed_
      -- CP-element group 404: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_324_Update/ca
      -- 
    ca_1196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_324_inst_ack_1, ack => access_T_CP_0_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	396 
    -- CP-element group 405: marked-predecessors 
    -- CP-element group 405: 	407 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	407 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_sample_start_
      -- CP-element group 405: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_Sample/rr
      -- 
    rr_1204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(405), ack => slice_328_inst_req_0); -- 
    access_T_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(396) & access_T_CP_0_elements(407);
      gj_access_T_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: marked-predecessors 
    -- CP-element group 406: 	432 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	408 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_update_start_
      -- CP-element group 406: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_Update/cr
      -- 
    cr_1209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(406), ack => slice_328_inst_req_1); -- 
    access_T_cp_element_group_406: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_406"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(432);
      gj_access_T_cp_element_group_406 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(406), clk => clk, reset => reset); --
    end block;
    -- CP-element group 407:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	405 
    -- CP-element group 407: successors 
    -- CP-element group 407: marked-successors 
    -- CP-element group 407: 	405 
    -- CP-element group 407: 	394 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_sample_completed_
      -- CP-element group 407: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_Sample/ra
      -- 
    ra_1205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_328_inst_ack_0, ack => access_T_CP_0_elements(407)); -- 
    -- CP-element group 408:  transition  input  bypass  pipeline-parent 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	406 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	431 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_update_completed_
      -- CP-element group 408: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_328_Update/ca
      -- 
    ca_1210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_328_inst_ack_1, ack => access_T_CP_0_elements(408)); -- 
    -- CP-element group 409:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	396 
    -- CP-element group 409: marked-predecessors 
    -- CP-element group 409: 	411 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	411 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_sample_start_
      -- CP-element group 409: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_Sample/$entry
      -- CP-element group 409: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_Sample/rr
      -- 
    rr_1218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(409), ack => slice_332_inst_req_0); -- 
    access_T_cp_element_group_409: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_409"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(396) & access_T_CP_0_elements(411);
      gj_access_T_cp_element_group_409 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(409), clk => clk, reset => reset); --
    end block;
    -- CP-element group 410:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: marked-predecessors 
    -- CP-element group 410: 	439 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	412 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_update_start_
      -- CP-element group 410: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_Update/cr
      -- 
    cr_1223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(410), ack => slice_332_inst_req_1); -- 
    access_T_cp_element_group_410: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_410"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(439);
      gj_access_T_cp_element_group_410 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(410), clk => clk, reset => reset); --
    end block;
    -- CP-element group 411:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	409 
    -- CP-element group 411: successors 
    -- CP-element group 411: marked-successors 
    -- CP-element group 411: 	409 
    -- CP-element group 411: 	394 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_sample_completed_
      -- CP-element group 411: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_Sample/$exit
      -- CP-element group 411: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_Sample/ra
      -- 
    ra_1219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_332_inst_ack_0, ack => access_T_CP_0_elements(411)); -- 
    -- CP-element group 412:  transition  input  bypass  pipeline-parent 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	410 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	438 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_update_completed_
      -- CP-element group 412: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_Update/$exit
      -- CP-element group 412: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_332_Update/ca
      -- 
    ca_1224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_332_inst_ack_1, ack => access_T_CP_0_elements(412)); -- 
    -- CP-element group 413:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	279 
    -- CP-element group 413: 	39 
    -- CP-element group 413: 	205 
    -- CP-element group 413: marked-predecessors 
    -- CP-element group 413: 	415 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	415 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_sample_start_
      -- CP-element group 413: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_Sample/$entry
      -- CP-element group 413: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_Sample/req
      -- 
    req_1232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(413), ack => W_send1_2_432_delayed_14_0_444_inst_req_0); -- 
    access_T_cp_element_group_413: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_413"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(279) & access_T_CP_0_elements(39) & access_T_CP_0_elements(205) & access_T_CP_0_elements(415);
      gj_access_T_cp_element_group_413 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(413), clk => clk, reset => reset); --
    end block;
    -- CP-element group 414:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: marked-predecessors 
    -- CP-element group 414: 	418 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	416 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_update_start_
      -- CP-element group 414: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_Update/req
      -- 
    req_1237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(414), ack => W_send1_2_432_delayed_14_0_444_inst_req_1); -- 
    access_T_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(418);
      gj_access_T_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	413 
    -- CP-element group 415: successors 
    -- CP-element group 415: marked-successors 
    -- CP-element group 415: 	277 
    -- CP-element group 415: 	201 
    -- CP-element group 415: 	35 
    -- CP-element group 415: 	413 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_sample_completed_
      -- CP-element group 415: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_Sample/ack
      -- 
    ack_1233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send1_2_432_delayed_14_0_444_inst_ack_0, ack => access_T_CP_0_elements(415)); -- 
    -- CP-element group 416:  transition  input  bypass  pipeline-parent 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	414 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_update_completed_
      -- CP-element group 416: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_446_Update/ack
      -- 
    ack_1238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send1_2_432_delayed_14_0_444_inst_ack_1, ack => access_T_CP_0_elements(416)); -- 
    -- CP-element group 417:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: 	400 
    -- CP-element group 417: marked-predecessors 
    -- CP-element group 417: 	440 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_sample_start_
      -- CP-element group 417: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_Sample/req
      -- 
    req_1246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(417), ack => WPIPE_input_pipe2_448_inst_req_0); -- 
    access_T_cp_element_group_417: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_417"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(416) & access_T_CP_0_elements(400) & access_T_CP_0_elements(440);
      gj_access_T_cp_element_group_417 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(417), clk => clk, reset => reset); --
    end block;
    -- CP-element group 418:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418: marked-successors 
    -- CP-element group 418: 	414 
    -- CP-element group 418: 	398 
    -- CP-element group 418:  members (6) 
      -- CP-element group 418: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_sample_completed_
      -- CP-element group 418: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_update_start_
      -- CP-element group 418: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_Sample/$exit
      -- CP-element group 418: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_Sample/ack
      -- CP-element group 418: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_Update/req
      -- 
    ack_1247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_448_inst_ack_0, ack => access_T_CP_0_elements(418)); -- 
    req_1251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(418), ack => WPIPE_input_pipe2_448_inst_req_1); -- 
    -- CP-element group 419:  transition  input  bypass  pipeline-parent 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	424 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_update_completed_
      -- CP-element group 419: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_Update/$exit
      -- CP-element group 419: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_448_Update/ack
      -- 
    ack_1252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_448_inst_ack_1, ack => access_T_CP_0_elements(419)); -- 
    -- CP-element group 420:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	279 
    -- CP-element group 420: 	39 
    -- CP-element group 420: 	205 
    -- CP-element group 420: 	123 
    -- CP-element group 420: marked-predecessors 
    -- CP-element group 420: 	422 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	422 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_sample_start_
      -- CP-element group 420: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_Sample/$entry
      -- CP-element group 420: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_Sample/req
      -- 
    req_1260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(420), ack => W_send2_2_436_delayed_14_0_451_inst_req_0); -- 
    access_T_cp_element_group_420: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_420"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(279) & access_T_CP_0_elements(39) & access_T_CP_0_elements(205) & access_T_CP_0_elements(123) & access_T_CP_0_elements(422);
      gj_access_T_cp_element_group_420 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(420), clk => clk, reset => reset); --
    end block;
    -- CP-element group 421:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: marked-predecessors 
    -- CP-element group 421: 	425 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	423 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_update_start_
      -- CP-element group 421: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_Update/$entry
      -- CP-element group 421: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_Update/req
      -- 
    req_1265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(421), ack => W_send2_2_436_delayed_14_0_451_inst_req_1); -- 
    access_T_cp_element_group_421: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_421"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(425);
      gj_access_T_cp_element_group_421 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(421), clk => clk, reset => reset); --
    end block;
    -- CP-element group 422:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	420 
    -- CP-element group 422: successors 
    -- CP-element group 422: marked-successors 
    -- CP-element group 422: 	277 
    -- CP-element group 422: 	201 
    -- CP-element group 422: 	35 
    -- CP-element group 422: 	420 
    -- CP-element group 422: 	119 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_sample_completed_
      -- CP-element group 422: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_Sample/$exit
      -- CP-element group 422: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_Sample/ack
      -- 
    ack_1261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send2_2_436_delayed_14_0_451_inst_ack_0, ack => access_T_CP_0_elements(422)); -- 
    -- CP-element group 423:  transition  input  bypass  pipeline-parent 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	421 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_update_completed_
      -- CP-element group 423: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_Update/$exit
      -- CP-element group 423: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_453_Update/ack
      -- 
    ack_1266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send2_2_436_delayed_14_0_451_inst_ack_1, ack => access_T_CP_0_elements(423)); -- 
    -- CP-element group 424:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	404 
    -- CP-element group 424: 	419 
    -- CP-element group 424: 	423 
    -- CP-element group 424: marked-predecessors 
    -- CP-element group 424: 	426 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_Sample/req
      -- 
    req_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(424), ack => WPIPE_input_pipe2_455_inst_req_0); -- 
    access_T_cp_element_group_424: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_424"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(404) & access_T_CP_0_elements(419) & access_T_CP_0_elements(423) & access_T_CP_0_elements(426);
      gj_access_T_cp_element_group_424 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(424), clk => clk, reset => reset); --
    end block;
    -- CP-element group 425:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425: marked-successors 
    -- CP-element group 425: 	421 
    -- CP-element group 425: 	402 
    -- CP-element group 425:  members (6) 
      -- CP-element group 425: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_sample_completed_
      -- CP-element group 425: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_update_start_
      -- CP-element group 425: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_Sample/ack
      -- CP-element group 425: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_Update/$entry
      -- CP-element group 425: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_Update/req
      -- 
    ack_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_455_inst_ack_0, ack => access_T_CP_0_elements(425)); -- 
    req_1279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(425), ack => WPIPE_input_pipe2_455_inst_req_1); -- 
    -- CP-element group 426:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	431 
    -- CP-element group 426: marked-successors 
    -- CP-element group 426: 	424 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_update_completed_
      -- CP-element group 426: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_455_Update/ack
      -- 
    ack_1280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_455_inst_ack_1, ack => access_T_CP_0_elements(426)); -- 
    -- CP-element group 427:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	279 
    -- CP-element group 427: 	39 
    -- CP-element group 427: 	205 
    -- CP-element group 427: 	123 
    -- CP-element group 427: marked-predecessors 
    -- CP-element group 427: 	429 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	429 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_Sample/req
      -- 
    req_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(427), ack => W_send3_2_440_delayed_14_0_458_inst_req_0); -- 
    access_T_cp_element_group_427: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_427"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(279) & access_T_CP_0_elements(39) & access_T_CP_0_elements(205) & access_T_CP_0_elements(123) & access_T_CP_0_elements(429);
      gj_access_T_cp_element_group_427 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(427), clk => clk, reset => reset); --
    end block;
    -- CP-element group 428:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: marked-predecessors 
    -- CP-element group 428: 	432 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	430 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_update_start_
      -- CP-element group 428: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_Update/$entry
      -- CP-element group 428: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_Update/req
      -- 
    req_1293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(428), ack => W_send3_2_440_delayed_14_0_458_inst_req_1); -- 
    access_T_cp_element_group_428: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_428"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(432);
      gj_access_T_cp_element_group_428 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(428), clk => clk, reset => reset); --
    end block;
    -- CP-element group 429:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	427 
    -- CP-element group 429: successors 
    -- CP-element group 429: marked-successors 
    -- CP-element group 429: 	277 
    -- CP-element group 429: 	201 
    -- CP-element group 429: 	35 
    -- CP-element group 429: 	427 
    -- CP-element group 429: 	119 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_sample_completed_
      -- CP-element group 429: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_Sample/$exit
      -- CP-element group 429: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_Sample/ack
      -- 
    ack_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send3_2_440_delayed_14_0_458_inst_ack_0, ack => access_T_CP_0_elements(429)); -- 
    -- CP-element group 430:  transition  input  bypass  pipeline-parent 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	428 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_update_completed_
      -- CP-element group 430: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_Update/$exit
      -- CP-element group 430: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_460_Update/ack
      -- 
    ack_1294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send3_2_440_delayed_14_0_458_inst_ack_1, ack => access_T_CP_0_elements(430)); -- 
    -- CP-element group 431:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	430 
    -- CP-element group 431: 	408 
    -- CP-element group 431: 	426 
    -- CP-element group 431: marked-predecessors 
    -- CP-element group 431: 	433 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	432 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_sample_start_
      -- CP-element group 431: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_Sample/$entry
      -- CP-element group 431: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_Sample/req
      -- 
    req_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(431), ack => WPIPE_input_pipe2_462_inst_req_0); -- 
    access_T_cp_element_group_431: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_431"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(430) & access_T_CP_0_elements(408) & access_T_CP_0_elements(426) & access_T_CP_0_elements(433);
      gj_access_T_cp_element_group_431 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(431), clk => clk, reset => reset); --
    end block;
    -- CP-element group 432:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	431 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432: marked-successors 
    -- CP-element group 432: 	406 
    -- CP-element group 432: 	428 
    -- CP-element group 432:  members (6) 
      -- CP-element group 432: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_update_start_
      -- CP-element group 432: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_Sample/ack
      -- CP-element group 432: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_Update/$entry
      -- CP-element group 432: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_Update/req
      -- 
    ack_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_462_inst_ack_0, ack => access_T_CP_0_elements(432)); -- 
    req_1307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(432), ack => WPIPE_input_pipe2_462_inst_req_1); -- 
    -- CP-element group 433:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	432 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	438 
    -- CP-element group 433: marked-successors 
    -- CP-element group 433: 	431 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_Update/$exit
      -- CP-element group 433: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_462_Update/ack
      -- 
    ack_1308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_462_inst_ack_1, ack => access_T_CP_0_elements(433)); -- 
    -- CP-element group 434:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	279 
    -- CP-element group 434: 	205 
    -- CP-element group 434: 	123 
    -- CP-element group 434: marked-predecessors 
    -- CP-element group 434: 	436 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	436 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_sample_start_
      -- CP-element group 434: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_Sample/$entry
      -- CP-element group 434: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_Sample/req
      -- 
    req_1316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(434), ack => W_send4_2_444_delayed_14_0_465_inst_req_0); -- 
    access_T_cp_element_group_434: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_434"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(279) & access_T_CP_0_elements(205) & access_T_CP_0_elements(123) & access_T_CP_0_elements(436);
      gj_access_T_cp_element_group_434 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(434), clk => clk, reset => reset); --
    end block;
    -- CP-element group 435:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: marked-predecessors 
    -- CP-element group 435: 	439 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	437 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_update_start_
      -- CP-element group 435: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_Update/$entry
      -- CP-element group 435: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_Update/req
      -- 
    req_1321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(435), ack => W_send4_2_444_delayed_14_0_465_inst_req_1); -- 
    access_T_cp_element_group_435: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_435"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(439);
      gj_access_T_cp_element_group_435 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(435), clk => clk, reset => reset); --
    end block;
    -- CP-element group 436:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	434 
    -- CP-element group 436: successors 
    -- CP-element group 436: marked-successors 
    -- CP-element group 436: 	277 
    -- CP-element group 436: 	201 
    -- CP-element group 436: 	434 
    -- CP-element group 436: 	119 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_sample_completed_
      -- CP-element group 436: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_Sample/$exit
      -- CP-element group 436: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_Sample/ack
      -- 
    ack_1317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send4_2_444_delayed_14_0_465_inst_ack_0, ack => access_T_CP_0_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass  pipeline-parent 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	435 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	438 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_update_completed_
      -- CP-element group 437: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_Update/$exit
      -- CP-element group 437: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_467_Update/ack
      -- 
    ack_1322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send4_2_444_delayed_14_0_465_inst_ack_1, ack => access_T_CP_0_elements(437)); -- 
    -- CP-element group 438:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	433 
    -- CP-element group 438: 	437 
    -- CP-element group 438: 	412 
    -- CP-element group 438: marked-predecessors 
    -- CP-element group 438: 	440 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	439 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_sample_start_
      -- CP-element group 438: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_Sample/$entry
      -- CP-element group 438: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_Sample/req
      -- 
    req_1330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(438), ack => WPIPE_input_pipe2_469_inst_req_0); -- 
    access_T_cp_element_group_438: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_438"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(433) & access_T_CP_0_elements(437) & access_T_CP_0_elements(412) & access_T_CP_0_elements(440);
      gj_access_T_cp_element_group_438 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(438), clk => clk, reset => reset); --
    end block;
    -- CP-element group 439:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	438 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439: marked-successors 
    -- CP-element group 439: 	435 
    -- CP-element group 439: 	410 
    -- CP-element group 439:  members (6) 
      -- CP-element group 439: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_sample_completed_
      -- CP-element group 439: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_update_start_
      -- CP-element group 439: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_Sample/$exit
      -- CP-element group 439: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_Sample/ack
      -- CP-element group 439: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_Update/$entry
      -- CP-element group 439: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_Update/req
      -- 
    ack_1331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_469_inst_ack_0, ack => access_T_CP_0_elements(439)); -- 
    req_1335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(439), ack => WPIPE_input_pipe2_469_inst_req_1); -- 
    -- CP-element group 440:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	552 
    -- CP-element group 440: marked-successors 
    -- CP-element group 440: 	438 
    -- CP-element group 440: 	417 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_update_completed_
      -- CP-element group 440: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_Update/$exit
      -- CP-element group 440: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_469_Update/ack
      -- 
    ack_1336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_469_inst_ack_1, ack => access_T_CP_0_elements(440)); -- 
    -- CP-element group 441:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	445 
    -- CP-element group 441: marked-predecessors 
    -- CP-element group 441: 	446 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	446 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_sample_start_
      -- CP-element group 441: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_request/$entry
      -- CP-element group 441: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_request/req
      -- 
    req_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(441), ack => addr_of_484_final_reg_req_0); -- 
    access_T_cp_element_group_441: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_441"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(445) & access_T_CP_0_elements(446);
      gj_access_T_cp_element_group_441 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(441), clk => clk, reset => reset); --
    end block;
    -- CP-element group 442:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	9 
    -- CP-element group 442: marked-predecessors 
    -- CP-element group 442: 	450 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	447 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_update_start_
      -- CP-element group 442: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_complete/$entry
      -- CP-element group 442: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_complete/req
      -- 
    req_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(442), ack => addr_of_484_final_reg_req_1); -- 
    access_T_cp_element_group_442: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_442"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(450);
      gj_access_T_cp_element_group_442 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(442), clk => clk, reset => reset); --
    end block;
    -- CP-element group 443:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	9 
    -- CP-element group 443: marked-predecessors 
    -- CP-element group 443: 	446 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	445 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_update_start
      -- CP-element group 443: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_Update/req
      -- 
    req_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(443), ack => array_obj_ref_483_index_offset_req_1); -- 
    access_T_cp_element_group_443: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_443"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(446);
      gj_access_T_cp_element_group_443 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(443), clk => clk, reset => reset); --
    end block;
    -- CP-element group 444:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	60 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	552 
    -- CP-element group 444: marked-successors 
    -- CP-element group 444: 	56 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_sample_complete
      -- CP-element group 444: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_Sample/ack
      -- 
    ack_1362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_483_index_offset_ack_0, ack => access_T_CP_0_elements(444)); -- 
    -- CP-element group 445:  transition  input  bypass  pipeline-parent 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	443 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	441 
    -- CP-element group 445:  members (8) 
      -- CP-element group 445: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_root_address_calculated
      -- CP-element group 445: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_offset_calculated
      -- CP-element group 445: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_final_index_sum_regn_Update/ack
      -- CP-element group 445: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_base_plus_offset/$entry
      -- CP-element group 445: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_base_plus_offset/$exit
      -- CP-element group 445: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_base_plus_offset/sum_rename_req
      -- CP-element group 445: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_483_base_plus_offset/sum_rename_ack
      -- 
    ack_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_483_index_offset_ack_1, ack => access_T_CP_0_elements(445)); -- 
    -- CP-element group 446:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	441 
    -- CP-element group 446: successors 
    -- CP-element group 446: marked-successors 
    -- CP-element group 446: 	441 
    -- CP-element group 446: 	443 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_sample_completed_
      -- CP-element group 446: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_request/$exit
      -- CP-element group 446: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_request/ack
      -- 
    ack_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_484_final_reg_ack_0, ack => access_T_CP_0_elements(446)); -- 
    -- CP-element group 447:  transition  input  bypass  pipeline-parent 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	442 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (19) 
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_plus_offset/sum_rename_req
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_word_addrgen/root_register_req
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_plus_offset/sum_rename_ack
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_word_addrgen/$entry
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_word_addrgen/root_register_ack
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_word_addrgen/$exit
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_plus_offset/$exit
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_plus_offset/$entry
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_addr_resize/base_resize_ack
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_addr_resize/base_resize_req
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_addr_resize/$exit
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_addr_resize/$entry
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_address_resized
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_root_address_calculated
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_update_completed_
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_complete/$exit
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_484_complete/ack
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_base_address_calculated
      -- CP-element group 447: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_word_address_calculated
      -- 
    ack_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_484_final_reg_ack_1, ack => access_T_CP_0_elements(447)); -- 
    -- CP-element group 448:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	447 
    -- CP-element group 448: marked-predecessors 
    -- CP-element group 448: 	450 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	450 
    -- CP-element group 448:  members (5) 
      -- CP-element group 448: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Sample/$entry
      -- CP-element group 448: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Sample/word_access_start/$entry
      -- CP-element group 448: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Sample/word_access_start/word_0/$entry
      -- CP-element group 448: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Sample/word_access_start/word_0/rr
      -- CP-element group 448: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_sample_start_
      -- 
    rr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(448), ack => ptr_deref_488_load_0_req_0); -- 
    access_T_cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(447) & access_T_CP_0_elements(450);
      gj_access_T_cp_element_group_448 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 449:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: marked-predecessors 
    -- CP-element group 449: 	454 
    -- CP-element group 449: 	458 
    -- CP-element group 449: 	462 
    -- CP-element group 449: 	466 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	451 
    -- CP-element group 449:  members (5) 
      -- CP-element group 449: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/word_access_complete/$entry
      -- CP-element group 449: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/word_access_complete/word_0/$entry
      -- CP-element group 449: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/word_access_complete/word_0/cr
      -- CP-element group 449: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_update_start_
      -- 
    cr_1426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(449), ack => ptr_deref_488_load_0_req_1); -- 
    access_T_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(454) & access_T_CP_0_elements(458) & access_T_CP_0_elements(462) & access_T_CP_0_elements(466);
      gj_access_T_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	448 
    -- CP-element group 450: successors 
    -- CP-element group 450: marked-successors 
    -- CP-element group 450: 	442 
    -- CP-element group 450: 	448 
    -- CP-element group 450:  members (5) 
      -- CP-element group 450: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Sample/word_access_start/$exit
      -- CP-element group 450: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Sample/word_access_start/word_0/$exit
      -- CP-element group 450: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Sample/$exit
      -- CP-element group 450: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Sample/word_access_start/word_0/ra
      -- CP-element group 450: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_sample_completed_
      -- 
    ra_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_488_load_0_ack_0, ack => access_T_CP_0_elements(450)); -- 
    -- CP-element group 451:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	449 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451: 	456 
    -- CP-element group 451: 	460 
    -- CP-element group 451: 	464 
    -- CP-element group 451:  members (9) 
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/word_access_complete/$exit
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/$exit
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/word_access_complete/word_0/$exit
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/ptr_deref_488_Merge/$entry
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/word_access_complete/word_0/ca
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/ptr_deref_488_Merge/$exit
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/ptr_deref_488_Merge/merge_req
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_Update/ptr_deref_488_Merge/merge_ack
      -- CP-element group 451: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_488_update_completed_
      -- 
    ca_1427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_488_load_0_ack_1, ack => access_T_CP_0_elements(451)); -- 
    -- CP-element group 452:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	451 
    -- CP-element group 452: marked-predecessors 
    -- CP-element group 452: 	454 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	454 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_Sample/$entry
      -- 
    rr_1440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(452), ack => slice_492_inst_req_0); -- 
    access_T_cp_element_group_452: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_452"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(451) & access_T_CP_0_elements(454);
      gj_access_T_cp_element_group_452 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(452), clk => clk, reset => reset); --
    end block;
    -- CP-element group 453:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: marked-predecessors 
    -- CP-element group 453: 	473 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	455 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_Update/$entry
      -- CP-element group 453: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_Update/cr
      -- CP-element group 453: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_update_start_
      -- 
    cr_1445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(453), ack => slice_492_inst_req_1); -- 
    access_T_cp_element_group_453: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_453"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(473);
      gj_access_T_cp_element_group_453 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(453), clk => clk, reset => reset); --
    end block;
    -- CP-element group 454:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	452 
    -- CP-element group 454: successors 
    -- CP-element group 454: marked-successors 
    -- CP-element group 454: 	449 
    -- CP-element group 454: 	452 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_sample_completed_
      -- CP-element group 454: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_Sample/$exit
      -- CP-element group 454: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_Sample/ra
      -- 
    ra_1441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_492_inst_ack_0, ack => access_T_CP_0_elements(454)); -- 
    -- CP-element group 455:  transition  input  bypass  pipeline-parent 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	453 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	472 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_Update/$exit
      -- CP-element group 455: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_Update/ca
      -- CP-element group 455: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_492_update_completed_
      -- 
    ca_1446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_492_inst_ack_1, ack => access_T_CP_0_elements(455)); -- 
    -- CP-element group 456:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	451 
    -- CP-element group 456: marked-predecessors 
    -- CP-element group 456: 	458 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	458 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_Sample/$entry
      -- CP-element group 456: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_sample_start_
      -- CP-element group 456: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_Sample/rr
      -- 
    rr_1454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(456), ack => slice_496_inst_req_0); -- 
    access_T_cp_element_group_456: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_456"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(451) & access_T_CP_0_elements(458);
      gj_access_T_cp_element_group_456 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(456), clk => clk, reset => reset); --
    end block;
    -- CP-element group 457:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: marked-predecessors 
    -- CP-element group 457: 	480 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	459 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_update_start_
      -- CP-element group 457: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_Update/cr
      -- CP-element group 457: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_Update/$entry
      -- 
    cr_1459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(457), ack => slice_496_inst_req_1); -- 
    access_T_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(480);
      gj_access_T_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	456 
    -- CP-element group 458: successors 
    -- CP-element group 458: marked-successors 
    -- CP-element group 458: 	449 
    -- CP-element group 458: 	456 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_sample_completed_
      -- CP-element group 458: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_Sample/ra
      -- CP-element group 458: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_Sample/$exit
      -- 
    ra_1455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_496_inst_ack_0, ack => access_T_CP_0_elements(458)); -- 
    -- CP-element group 459:  transition  input  bypass  pipeline-parent 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	457 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	479 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_update_completed_
      -- CP-element group 459: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_Update/ca
      -- CP-element group 459: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_496_Update/$exit
      -- 
    ca_1460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_496_inst_ack_1, ack => access_T_CP_0_elements(459)); -- 
    -- CP-element group 460:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	451 
    -- CP-element group 460: marked-predecessors 
    -- CP-element group 460: 	462 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	462 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_Sample/rr
      -- CP-element group 460: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_sample_start_
      -- 
    rr_1468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(460), ack => slice_500_inst_req_0); -- 
    access_T_cp_element_group_460: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_460"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(451) & access_T_CP_0_elements(462);
      gj_access_T_cp_element_group_460 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(460), clk => clk, reset => reset); --
    end block;
    -- CP-element group 461:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: marked-predecessors 
    -- CP-element group 461: 	487 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	463 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_update_start_
      -- 
    cr_1473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(461), ack => slice_500_inst_req_1); -- 
    access_T_cp_element_group_461: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_461"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(487);
      gj_access_T_cp_element_group_461 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(461), clk => clk, reset => reset); --
    end block;
    -- CP-element group 462:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	460 
    -- CP-element group 462: successors 
    -- CP-element group 462: marked-successors 
    -- CP-element group 462: 	449 
    -- CP-element group 462: 	460 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_Sample/ra
      -- CP-element group 462: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_Sample/$exit
      -- CP-element group 462: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_sample_completed_
      -- 
    ra_1469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_500_inst_ack_0, ack => access_T_CP_0_elements(462)); -- 
    -- CP-element group 463:  transition  input  bypass  pipeline-parent 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	461 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	486 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_Update/ca
      -- CP-element group 463: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_Update/$exit
      -- CP-element group 463: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_500_update_completed_
      -- 
    ca_1474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_500_inst_ack_1, ack => access_T_CP_0_elements(463)); -- 
    -- CP-element group 464:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	451 
    -- CP-element group 464: marked-predecessors 
    -- CP-element group 464: 	466 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	466 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_Sample/rr
      -- CP-element group 464: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_Sample/$entry
      -- CP-element group 464: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_sample_start_
      -- 
    rr_1482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(464), ack => slice_504_inst_req_0); -- 
    access_T_cp_element_group_464: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_464"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(451) & access_T_CP_0_elements(466);
      gj_access_T_cp_element_group_464 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(464), clk => clk, reset => reset); --
    end block;
    -- CP-element group 465:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: marked-predecessors 
    -- CP-element group 465: 	494 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	467 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_Update/cr
      -- CP-element group 465: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_update_start_
      -- CP-element group 465: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_Update/$entry
      -- 
    cr_1487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(465), ack => slice_504_inst_req_1); -- 
    access_T_cp_element_group_465: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_465"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(494);
      gj_access_T_cp_element_group_465 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(465), clk => clk, reset => reset); --
    end block;
    -- CP-element group 466:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	464 
    -- CP-element group 466: successors 
    -- CP-element group 466: marked-successors 
    -- CP-element group 466: 	449 
    -- CP-element group 466: 	464 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_Sample/$exit
      -- CP-element group 466: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_Sample/ra
      -- CP-element group 466: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_sample_completed_
      -- 
    ra_1483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_504_inst_ack_0, ack => access_T_CP_0_elements(466)); -- 
    -- CP-element group 467:  transition  input  bypass  pipeline-parent 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	465 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	493 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_update_completed_
      -- CP-element group 467: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_Update/ca
      -- CP-element group 467: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_504_Update/$exit
      -- 
    ca_1488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_504_inst_ack_1, ack => access_T_CP_0_elements(467)); -- 
    -- CP-element group 468:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	298 
    -- CP-element group 468: 	60 
    -- CP-element group 468: 	224 
    -- CP-element group 468: marked-predecessors 
    -- CP-element group 468: 	470 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	470 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_Sample/req
      -- CP-element group 468: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_sample_start_
      -- CP-element group 468: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_Sample/$entry
      -- 
    req_1496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(468), ack => W_send1_3_592_delayed_14_0_616_inst_req_0); -- 
    access_T_cp_element_group_468: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_468"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(298) & access_T_CP_0_elements(60) & access_T_CP_0_elements(224) & access_T_CP_0_elements(470);
      gj_access_T_cp_element_group_468 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(468), clk => clk, reset => reset); --
    end block;
    -- CP-element group 469:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: marked-predecessors 
    -- CP-element group 469: 	473 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	471 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_update_start_
      -- CP-element group 469: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_Update/req
      -- 
    req_1501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(469), ack => W_send1_3_592_delayed_14_0_616_inst_req_1); -- 
    access_T_cp_element_group_469: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_469"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(473);
      gj_access_T_cp_element_group_469 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(469), clk => clk, reset => reset); --
    end block;
    -- CP-element group 470:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	468 
    -- CP-element group 470: successors 
    -- CP-element group 470: marked-successors 
    -- CP-element group 470: 	294 
    -- CP-element group 470: 	56 
    -- CP-element group 470: 	220 
    -- CP-element group 470: 	468 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_Sample/ack
      -- CP-element group 470: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_Sample/$exit
      -- CP-element group 470: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_sample_completed_
      -- 
    ack_1497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send1_3_592_delayed_14_0_616_inst_ack_0, ack => access_T_CP_0_elements(470)); -- 
    -- CP-element group 471:  transition  input  bypass  pipeline-parent 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	469 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	472 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_update_completed_
      -- CP-element group 471: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_Update/$exit
      -- CP-element group 471: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_618_Update/ack
      -- 
    ack_1502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send1_3_592_delayed_14_0_616_inst_ack_1, ack => access_T_CP_0_elements(471)); -- 
    -- CP-element group 472:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	471 
    -- CP-element group 472: 	455 
    -- CP-element group 472: marked-predecessors 
    -- CP-element group 472: 	495 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_Sample/req
      -- 
    req_1510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(472), ack => WPIPE_input_pipe3_620_inst_req_0); -- 
    access_T_cp_element_group_472: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_472"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(471) & access_T_CP_0_elements(455) & access_T_CP_0_elements(495);
      gj_access_T_cp_element_group_472 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(472), clk => clk, reset => reset); --
    end block;
    -- CP-element group 473:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473: marked-successors 
    -- CP-element group 473: 	469 
    -- CP-element group 473: 	453 
    -- CP-element group 473:  members (6) 
      -- CP-element group 473: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_update_start_
      -- CP-element group 473: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_sample_completed_
      -- CP-element group 473: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_Sample/$exit
      -- CP-element group 473: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_Sample/ack
      -- CP-element group 473: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_Update/$entry
      -- CP-element group 473: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_Update/req
      -- 
    ack_1511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_620_inst_ack_0, ack => access_T_CP_0_elements(473)); -- 
    req_1515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(473), ack => WPIPE_input_pipe3_620_inst_req_1); -- 
    -- CP-element group 474:  transition  input  bypass  pipeline-parent 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	479 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_update_completed_
      -- CP-element group 474: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_Update/$exit
      -- CP-element group 474: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_620_Update/ack
      -- 
    ack_1516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_620_inst_ack_1, ack => access_T_CP_0_elements(474)); -- 
    -- CP-element group 475:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	144 
    -- CP-element group 475: 	298 
    -- CP-element group 475: 	60 
    -- CP-element group 475: 	224 
    -- CP-element group 475: marked-predecessors 
    -- CP-element group 475: 	477 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	477 
    -- CP-element group 475:  members (3) 
      -- CP-element group 475: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_Sample/req
      -- CP-element group 475: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_Sample/$entry
      -- 
    req_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(475), ack => W_send2_3_596_delayed_14_0_623_inst_req_0); -- 
    access_T_cp_element_group_475: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_475"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(144) & access_T_CP_0_elements(298) & access_T_CP_0_elements(60) & access_T_CP_0_elements(224) & access_T_CP_0_elements(477);
      gj_access_T_cp_element_group_475 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(475), clk => clk, reset => reset); --
    end block;
    -- CP-element group 476:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: marked-predecessors 
    -- CP-element group 476: 	480 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	478 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_update_start_
      -- CP-element group 476: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_Update/req
      -- CP-element group 476: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_Update/$entry
      -- 
    req_1529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(476), ack => W_send2_3_596_delayed_14_0_623_inst_req_1); -- 
    access_T_cp_element_group_476: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_476"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(480);
      gj_access_T_cp_element_group_476 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(476), clk => clk, reset => reset); --
    end block;
    -- CP-element group 477:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	475 
    -- CP-element group 477: successors 
    -- CP-element group 477: marked-successors 
    -- CP-element group 477: 	140 
    -- CP-element group 477: 	294 
    -- CP-element group 477: 	56 
    -- CP-element group 477: 	475 
    -- CP-element group 477: 	220 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_sample_completed_
      -- CP-element group 477: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_Sample/ack
      -- CP-element group 477: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_Sample/$exit
      -- 
    ack_1525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send2_3_596_delayed_14_0_623_inst_ack_0, ack => access_T_CP_0_elements(477)); -- 
    -- CP-element group 478:  transition  input  bypass  pipeline-parent 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	476 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	479 
    -- CP-element group 478:  members (3) 
      -- CP-element group 478: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_Update/ack
      -- CP-element group 478: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_Update/$exit
      -- CP-element group 478: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_625_update_completed_
      -- 
    ack_1530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send2_3_596_delayed_14_0_623_inst_ack_1, ack => access_T_CP_0_elements(478)); -- 
    -- CP-element group 479:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	474 
    -- CP-element group 479: 	478 
    -- CP-element group 479: 	459 
    -- CP-element group 479: marked-predecessors 
    -- CP-element group 479: 	481 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_sample_start_
      -- CP-element group 479: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_Sample/$entry
      -- CP-element group 479: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_Sample/req
      -- 
    req_1538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(479), ack => WPIPE_input_pipe3_627_inst_req_0); -- 
    access_T_cp_element_group_479: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_479"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(474) & access_T_CP_0_elements(478) & access_T_CP_0_elements(459) & access_T_CP_0_elements(481);
      gj_access_T_cp_element_group_479 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(479), clk => clk, reset => reset); --
    end block;
    -- CP-element group 480:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480: marked-successors 
    -- CP-element group 480: 	476 
    -- CP-element group 480: 	457 
    -- CP-element group 480:  members (6) 
      -- CP-element group 480: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_sample_completed_
      -- CP-element group 480: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_update_start_
      -- CP-element group 480: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_Sample/$exit
      -- CP-element group 480: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_Update/req
      -- CP-element group 480: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_Sample/ack
      -- CP-element group 480: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_Update/$entry
      -- 
    ack_1539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_627_inst_ack_0, ack => access_T_CP_0_elements(480)); -- 
    req_1543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(480), ack => WPIPE_input_pipe3_627_inst_req_1); -- 
    -- CP-element group 481:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	486 
    -- CP-element group 481: marked-successors 
    -- CP-element group 481: 	479 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_update_completed_
      -- CP-element group 481: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_Update/$exit
      -- CP-element group 481: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_627_Update/ack
      -- 
    ack_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_627_inst_ack_1, ack => access_T_CP_0_elements(481)); -- 
    -- CP-element group 482:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	144 
    -- CP-element group 482: 	298 
    -- CP-element group 482: 	60 
    -- CP-element group 482: 	224 
    -- CP-element group 482: marked-predecessors 
    -- CP-element group 482: 	484 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	484 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_Sample/req
      -- CP-element group 482: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_sample_start_
      -- 
    req_1552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(482), ack => W_send3_3_600_delayed_14_0_630_inst_req_0); -- 
    access_T_cp_element_group_482: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_482"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(144) & access_T_CP_0_elements(298) & access_T_CP_0_elements(60) & access_T_CP_0_elements(224) & access_T_CP_0_elements(484);
      gj_access_T_cp_element_group_482 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(482), clk => clk, reset => reset); --
    end block;
    -- CP-element group 483:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: marked-predecessors 
    -- CP-element group 483: 	487 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	485 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_Update/req
      -- CP-element group 483: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_update_start_
      -- 
    req_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(483), ack => W_send3_3_600_delayed_14_0_630_inst_req_1); -- 
    access_T_cp_element_group_483: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_483"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(487);
      gj_access_T_cp_element_group_483 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(483), clk => clk, reset => reset); --
    end block;
    -- CP-element group 484:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	482 
    -- CP-element group 484: successors 
    -- CP-element group 484: marked-successors 
    -- CP-element group 484: 	140 
    -- CP-element group 484: 	294 
    -- CP-element group 484: 	56 
    -- CP-element group 484: 	482 
    -- CP-element group 484: 	220 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_Sample/ack
      -- CP-element group 484: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_sample_completed_
      -- 
    ack_1553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send3_3_600_delayed_14_0_630_inst_ack_0, ack => access_T_CP_0_elements(484)); -- 
    -- CP-element group 485:  transition  input  bypass  pipeline-parent 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	483 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	486 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_Update/ack
      -- CP-element group 485: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_632_update_completed_
      -- 
    ack_1558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send3_3_600_delayed_14_0_630_inst_ack_1, ack => access_T_CP_0_elements(485)); -- 
    -- CP-element group 486:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	481 
    -- CP-element group 486: 	485 
    -- CP-element group 486: 	463 
    -- CP-element group 486: marked-predecessors 
    -- CP-element group 486: 	488 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_Sample/req
      -- CP-element group 486: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_sample_start_
      -- 
    req_1566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(486), ack => WPIPE_input_pipe3_634_inst_req_0); -- 
    access_T_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(481) & access_T_CP_0_elements(485) & access_T_CP_0_elements(463) & access_T_CP_0_elements(488);
      gj_access_T_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487: marked-successors 
    -- CP-element group 487: 	483 
    -- CP-element group 487: 	461 
    -- CP-element group 487:  members (6) 
      -- CP-element group 487: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_Update/req
      -- CP-element group 487: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_Update/$entry
      -- CP-element group 487: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_Sample/ack
      -- CP-element group 487: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_Sample/$exit
      -- CP-element group 487: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_update_start_
      -- CP-element group 487: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_sample_completed_
      -- 
    ack_1567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_634_inst_ack_0, ack => access_T_CP_0_elements(487)); -- 
    req_1571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(487), ack => WPIPE_input_pipe3_634_inst_req_1); -- 
    -- CP-element group 488:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	493 
    -- CP-element group 488: marked-successors 
    -- CP-element group 488: 	486 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_Update/ack
      -- CP-element group 488: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_Update/$exit
      -- CP-element group 488: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_634_update_completed_
      -- 
    ack_1572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_634_inst_ack_1, ack => access_T_CP_0_elements(488)); -- 
    -- CP-element group 489:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	144 
    -- CP-element group 489: 	298 
    -- CP-element group 489: 	224 
    -- CP-element group 489: marked-predecessors 
    -- CP-element group 489: 	491 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	491 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_Sample/req
      -- 
    req_1580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(489), ack => W_send4_3_604_delayed_14_0_637_inst_req_0); -- 
    access_T_cp_element_group_489: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_489"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(144) & access_T_CP_0_elements(298) & access_T_CP_0_elements(224) & access_T_CP_0_elements(491);
      gj_access_T_cp_element_group_489 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(489), clk => clk, reset => reset); --
    end block;
    -- CP-element group 490:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: marked-predecessors 
    -- CP-element group 490: 	494 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	492 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_update_start_
      -- CP-element group 490: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_Update/req
      -- CP-element group 490: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_Update/$entry
      -- 
    req_1585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(490), ack => W_send4_3_604_delayed_14_0_637_inst_req_1); -- 
    access_T_cp_element_group_490: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_490"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(494);
      gj_access_T_cp_element_group_490 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(490), clk => clk, reset => reset); --
    end block;
    -- CP-element group 491:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	489 
    -- CP-element group 491: successors 
    -- CP-element group 491: marked-successors 
    -- CP-element group 491: 	140 
    -- CP-element group 491: 	294 
    -- CP-element group 491: 	489 
    -- CP-element group 491: 	220 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_sample_completed_
      -- CP-element group 491: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_Sample/ack
      -- 
    ack_1581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send4_3_604_delayed_14_0_637_inst_ack_0, ack => access_T_CP_0_elements(491)); -- 
    -- CP-element group 492:  transition  input  bypass  pipeline-parent 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	490 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492:  members (3) 
      -- CP-element group 492: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_update_completed_
      -- CP-element group 492: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_639_Update/ack
      -- 
    ack_1586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send4_3_604_delayed_14_0_637_inst_ack_1, ack => access_T_CP_0_elements(492)); -- 
    -- CP-element group 493:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	488 
    -- CP-element group 493: 	492 
    -- CP-element group 493: 	467 
    -- CP-element group 493: marked-predecessors 
    -- CP-element group 493: 	495 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_sample_start_
      -- CP-element group 493: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_Sample/$entry
      -- CP-element group 493: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_Sample/req
      -- 
    req_1594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(493), ack => WPIPE_input_pipe3_641_inst_req_0); -- 
    access_T_cp_element_group_493: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_493"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(488) & access_T_CP_0_elements(492) & access_T_CP_0_elements(467) & access_T_CP_0_elements(495);
      gj_access_T_cp_element_group_493 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(493), clk => clk, reset => reset); --
    end block;
    -- CP-element group 494:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	493 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494: marked-successors 
    -- CP-element group 494: 	490 
    -- CP-element group 494: 	465 
    -- CP-element group 494:  members (6) 
      -- CP-element group 494: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_sample_completed_
      -- CP-element group 494: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_update_start_
      -- CP-element group 494: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_Sample/$exit
      -- CP-element group 494: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_Sample/ack
      -- CP-element group 494: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_Update/$entry
      -- CP-element group 494: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_Update/req
      -- 
    ack_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_641_inst_ack_0, ack => access_T_CP_0_elements(494)); -- 
    req_1599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(494), ack => WPIPE_input_pipe3_641_inst_req_1); -- 
    -- CP-element group 495:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	552 
    -- CP-element group 495: marked-successors 
    -- CP-element group 495: 	472 
    -- CP-element group 495: 	493 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_update_completed_
      -- CP-element group 495: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_Update/$exit
      -- CP-element group 495: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_641_Update/ack
      -- 
    ack_1600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_641_inst_ack_1, ack => access_T_CP_0_elements(495)); -- 
    -- CP-element group 496:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	500 
    -- CP-element group 496: marked-predecessors 
    -- CP-element group 496: 	501 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	501 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_sample_start_
      -- CP-element group 496: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_request/req
      -- CP-element group 496: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_request/$entry
      -- 
    req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(496), ack => addr_of_656_final_reg_req_0); -- 
    access_T_cp_element_group_496: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_496"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(500) & access_T_CP_0_elements(501);
      gj_access_T_cp_element_group_496 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(496), clk => clk, reset => reset); --
    end block;
    -- CP-element group 497:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	9 
    -- CP-element group 497: marked-predecessors 
    -- CP-element group 497: 	505 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	502 
    -- CP-element group 497:  members (3) 
      -- CP-element group 497: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_update_start_
      -- CP-element group 497: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_complete/req
      -- CP-element group 497: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_complete/$entry
      -- 
    req_1645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(497), ack => addr_of_656_final_reg_req_1); -- 
    access_T_cp_element_group_497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(505);
      gj_access_T_cp_element_group_497 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 498:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	9 
    -- CP-element group 498: marked-predecessors 
    -- CP-element group 498: 	501 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	500 
    -- CP-element group 498:  members (3) 
      -- CP-element group 498: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_Update/req
      -- CP-element group 498: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_update_start
      -- 
    req_1630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(498), ack => array_obj_ref_655_index_offset_req_1); -- 
    access_T_cp_element_group_498: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_498"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(501);
      gj_access_T_cp_element_group_498 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(498), clk => clk, reset => reset); --
    end block;
    -- CP-element group 499:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	81 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	552 
    -- CP-element group 499: marked-successors 
    -- CP-element group 499: 	77 
    -- CP-element group 499:  members (3) 
      -- CP-element group 499: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_sample_complete
      -- CP-element group 499: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_Sample/$exit
      -- CP-element group 499: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_Sample/ack
      -- 
    ack_1626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_655_index_offset_ack_0, ack => access_T_CP_0_elements(499)); -- 
    -- CP-element group 500:  transition  input  bypass  pipeline-parent 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	498 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	496 
    -- CP-element group 500:  members (8) 
      -- CP-element group 500: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_Update/$exit
      -- CP-element group 500: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_final_index_sum_regn_Update/ack
      -- CP-element group 500: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_base_plus_offset/sum_rename_ack
      -- CP-element group 500: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_base_plus_offset/sum_rename_req
      -- CP-element group 500: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_base_plus_offset/$exit
      -- CP-element group 500: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_base_plus_offset/$entry
      -- CP-element group 500: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_offset_calculated
      -- CP-element group 500: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_655_root_address_calculated
      -- 
    ack_1631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_655_index_offset_ack_1, ack => access_T_CP_0_elements(500)); -- 
    -- CP-element group 501:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	496 
    -- CP-element group 501: successors 
    -- CP-element group 501: marked-successors 
    -- CP-element group 501: 	496 
    -- CP-element group 501: 	498 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_sample_completed_
      -- CP-element group 501: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_request/ack
      -- CP-element group 501: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_request/$exit
      -- 
    ack_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_656_final_reg_ack_0, ack => access_T_CP_0_elements(501)); -- 
    -- CP-element group 502:  transition  input  bypass  pipeline-parent 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	497 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	503 
    -- CP-element group 502:  members (19) 
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_addr_resize/base_resize_req
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_addr_resize/base_resize_ack
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_addr_resize/$entry
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_address_calculated
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_word_address_calculated
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_plus_offset/$entry
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_root_address_calculated
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_address_resized
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_word_addrgen/root_register_ack
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_complete/ack
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_complete/$exit
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_addr_resize/$exit
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_word_addrgen/root_register_req
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_word_addrgen/$exit
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_word_addrgen/$entry
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_plus_offset/sum_rename_ack
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_plus_offset/sum_rename_req
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_base_plus_offset/$exit
      -- CP-element group 502: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_656_update_completed_
      -- 
    ack_1646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_656_final_reg_ack_1, ack => access_T_CP_0_elements(502)); -- 
    -- CP-element group 503:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	502 
    -- CP-element group 503: marked-predecessors 
    -- CP-element group 503: 	505 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	505 
    -- CP-element group 503:  members (5) 
      -- CP-element group 503: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_sample_start_
      -- CP-element group 503: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Sample/word_access_start/$entry
      -- CP-element group 503: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Sample/word_access_start/word_0/$entry
      -- CP-element group 503: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Sample/word_access_start/word_0/rr
      -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(503), ack => ptr_deref_660_load_0_req_0); -- 
    access_T_cp_element_group_503: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_503"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(502) & access_T_CP_0_elements(505);
      gj_access_T_cp_element_group_503 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(503), clk => clk, reset => reset); --
    end block;
    -- CP-element group 504:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: marked-predecessors 
    -- CP-element group 504: 	509 
    -- CP-element group 504: 	513 
    -- CP-element group 504: 	517 
    -- CP-element group 504: 	521 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	506 
    -- CP-element group 504:  members (5) 
      -- CP-element group 504: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_update_start_
      -- CP-element group 504: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/word_access_complete/word_0/cr
      -- CP-element group 504: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/word_access_complete/word_0/$entry
      -- CP-element group 504: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/word_access_complete/$entry
      -- CP-element group 504: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/$entry
      -- 
    cr_1690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(504), ack => ptr_deref_660_load_0_req_1); -- 
    access_T_cp_element_group_504: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_504"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(509) & access_T_CP_0_elements(513) & access_T_CP_0_elements(517) & access_T_CP_0_elements(521);
      gj_access_T_cp_element_group_504 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(504), clk => clk, reset => reset); --
    end block;
    -- CP-element group 505:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	503 
    -- CP-element group 505: successors 
    -- CP-element group 505: marked-successors 
    -- CP-element group 505: 	497 
    -- CP-element group 505: 	503 
    -- CP-element group 505:  members (5) 
      -- CP-element group 505: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Sample/$exit
      -- CP-element group 505: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_sample_completed_
      -- CP-element group 505: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Sample/word_access_start/word_0/$exit
      -- CP-element group 505: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Sample/word_access_start/$exit
      -- CP-element group 505: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Sample/word_access_start/word_0/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_660_load_0_ack_0, ack => access_T_CP_0_elements(505)); -- 
    -- CP-element group 506:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	504 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	507 
    -- CP-element group 506: 	511 
    -- CP-element group 506: 	515 
    -- CP-element group 506: 	519 
    -- CP-element group 506:  members (9) 
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_update_completed_
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/ptr_deref_660_Merge/merge_ack
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/ptr_deref_660_Merge/merge_req
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/ptr_deref_660_Merge/$exit
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/ptr_deref_660_Merge/$entry
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/word_access_complete/word_0/ca
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/word_access_complete/word_0/$exit
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/word_access_complete/$exit
      -- CP-element group 506: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_660_Update/$exit
      -- 
    ca_1691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_660_load_0_ack_1, ack => access_T_CP_0_elements(506)); -- 
    -- CP-element group 507:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	506 
    -- CP-element group 507: marked-predecessors 
    -- CP-element group 507: 	509 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	509 
    -- CP-element group 507:  members (3) 
      -- CP-element group 507: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_Sample/rr
      -- 
    rr_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(507), ack => slice_664_inst_req_0); -- 
    access_T_cp_element_group_507: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_507"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(506) & access_T_CP_0_elements(509);
      gj_access_T_cp_element_group_507 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(507), clk => clk, reset => reset); --
    end block;
    -- CP-element group 508:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: marked-predecessors 
    -- CP-element group 508: 	528 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	510 
    -- CP-element group 508:  members (3) 
      -- CP-element group 508: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_Update/cr
      -- CP-element group 508: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_Update/$entry
      -- CP-element group 508: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_update_start_
      -- 
    cr_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(508), ack => slice_664_inst_req_1); -- 
    access_T_cp_element_group_508: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_508"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(528);
      gj_access_T_cp_element_group_508 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(508), clk => clk, reset => reset); --
    end block;
    -- CP-element group 509:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	507 
    -- CP-element group 509: successors 
    -- CP-element group 509: marked-successors 
    -- CP-element group 509: 	504 
    -- CP-element group 509: 	507 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_sample_completed_
      -- CP-element group 509: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_Sample/$exit
      -- CP-element group 509: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_Sample/ra
      -- 
    ra_1705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_664_inst_ack_0, ack => access_T_CP_0_elements(509)); -- 
    -- CP-element group 510:  transition  input  bypass  pipeline-parent 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	508 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	527 
    -- CP-element group 510:  members (3) 
      -- CP-element group 510: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_Update/$exit
      -- CP-element group 510: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_Update/ca
      -- CP-element group 510: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_664_update_completed_
      -- 
    ca_1710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_664_inst_ack_1, ack => access_T_CP_0_elements(510)); -- 
    -- CP-element group 511:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	506 
    -- CP-element group 511: marked-predecessors 
    -- CP-element group 511: 	513 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	513 
    -- CP-element group 511:  members (3) 
      -- CP-element group 511: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_sample_start_
      -- CP-element group 511: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_Sample/rr
      -- CP-element group 511: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_Sample/$entry
      -- 
    rr_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(511), ack => slice_668_inst_req_0); -- 
    access_T_cp_element_group_511: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_511"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(506) & access_T_CP_0_elements(513);
      gj_access_T_cp_element_group_511 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(511), clk => clk, reset => reset); --
    end block;
    -- CP-element group 512:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: marked-predecessors 
    -- CP-element group 512: 	535 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	514 
    -- CP-element group 512:  members (3) 
      -- CP-element group 512: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_Update/cr
      -- CP-element group 512: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_Update/$entry
      -- CP-element group 512: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_update_start_
      -- 
    cr_1723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(512), ack => slice_668_inst_req_1); -- 
    access_T_cp_element_group_512: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_512"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(535);
      gj_access_T_cp_element_group_512 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(512), clk => clk, reset => reset); --
    end block;
    -- CP-element group 513:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	511 
    -- CP-element group 513: successors 
    -- CP-element group 513: marked-successors 
    -- CP-element group 513: 	504 
    -- CP-element group 513: 	511 
    -- CP-element group 513:  members (3) 
      -- CP-element group 513: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_sample_completed_
      -- CP-element group 513: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_Sample/ra
      -- CP-element group 513: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_Sample/$exit
      -- 
    ra_1719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_668_inst_ack_0, ack => access_T_CP_0_elements(513)); -- 
    -- CP-element group 514:  transition  input  bypass  pipeline-parent 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	512 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	534 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_Update/$exit
      -- CP-element group 514: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_Update/ca
      -- CP-element group 514: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_668_update_completed_
      -- 
    ca_1724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_668_inst_ack_1, ack => access_T_CP_0_elements(514)); -- 
    -- CP-element group 515:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	506 
    -- CP-element group 515: marked-predecessors 
    -- CP-element group 515: 	517 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	517 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_Sample/$entry
      -- CP-element group 515: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_Sample/rr
      -- CP-element group 515: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_sample_start_
      -- 
    rr_1732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(515), ack => slice_672_inst_req_0); -- 
    access_T_cp_element_group_515: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_515"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(506) & access_T_CP_0_elements(517);
      gj_access_T_cp_element_group_515 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(515), clk => clk, reset => reset); --
    end block;
    -- CP-element group 516:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: marked-predecessors 
    -- CP-element group 516: 	542 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	518 
    -- CP-element group 516:  members (3) 
      -- CP-element group 516: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_Update/$entry
      -- CP-element group 516: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_update_start_
      -- CP-element group 516: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_Update/cr
      -- 
    cr_1737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(516), ack => slice_672_inst_req_1); -- 
    access_T_cp_element_group_516: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_516"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(542);
      gj_access_T_cp_element_group_516 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(516), clk => clk, reset => reset); --
    end block;
    -- CP-element group 517:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	515 
    -- CP-element group 517: successors 
    -- CP-element group 517: marked-successors 
    -- CP-element group 517: 	504 
    -- CP-element group 517: 	515 
    -- CP-element group 517:  members (3) 
      -- CP-element group 517: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_Sample/ra
      -- CP-element group 517: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_Sample/$exit
      -- CP-element group 517: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_sample_completed_
      -- 
    ra_1733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_672_inst_ack_0, ack => access_T_CP_0_elements(517)); -- 
    -- CP-element group 518:  transition  input  bypass  pipeline-parent 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	516 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	541 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_update_completed_
      -- CP-element group 518: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_Update/ca
      -- CP-element group 518: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_672_Update/$exit
      -- 
    ca_1738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_672_inst_ack_1, ack => access_T_CP_0_elements(518)); -- 
    -- CP-element group 519:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	506 
    -- CP-element group 519: marked-predecessors 
    -- CP-element group 519: 	521 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	521 
    -- CP-element group 519:  members (3) 
      -- CP-element group 519: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_Sample/$entry
      -- CP-element group 519: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_sample_start_
      -- CP-element group 519: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_Sample/rr
      -- 
    rr_1746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(519), ack => slice_676_inst_req_0); -- 
    access_T_cp_element_group_519: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_519"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(506) & access_T_CP_0_elements(521);
      gj_access_T_cp_element_group_519 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(519), clk => clk, reset => reset); --
    end block;
    -- CP-element group 520:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: marked-predecessors 
    -- CP-element group 520: 	549 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	522 
    -- CP-element group 520:  members (3) 
      -- CP-element group 520: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_update_start_
      -- CP-element group 520: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_Update/$entry
      -- 
    cr_1751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(520), ack => slice_676_inst_req_1); -- 
    access_T_cp_element_group_520: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_520"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(549);
      gj_access_T_cp_element_group_520 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(520), clk => clk, reset => reset); --
    end block;
    -- CP-element group 521:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	519 
    -- CP-element group 521: successors 
    -- CP-element group 521: marked-successors 
    -- CP-element group 521: 	504 
    -- CP-element group 521: 	519 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_Sample/$exit
      -- CP-element group 521: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_sample_completed_
      -- CP-element group 521: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_Sample/ra
      -- 
    ra_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_676_inst_ack_0, ack => access_T_CP_0_elements(521)); -- 
    -- CP-element group 522:  transition  input  bypass  pipeline-parent 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	520 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	548 
    -- CP-element group 522:  members (3) 
      -- CP-element group 522: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_Update/ca
      -- CP-element group 522: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_update_completed_
      -- CP-element group 522: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/slice_676_Update/$exit
      -- 
    ca_1752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 522_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_676_inst_ack_1, ack => access_T_CP_0_elements(522)); -- 
    -- CP-element group 523:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	317 
    -- CP-element group 523: 	81 
    -- CP-element group 523: 	243 
    -- CP-element group 523: marked-predecessors 
    -- CP-element group 523: 	525 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	525 
    -- CP-element group 523:  members (3) 
      -- CP-element group 523: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_Sample/req
      -- CP-element group 523: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_Sample/$entry
      -- CP-element group 523: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_sample_start_
      -- 
    req_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(523), ack => W_send1_4_752_delayed_14_0_788_inst_req_0); -- 
    access_T_cp_element_group_523: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_523"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(317) & access_T_CP_0_elements(81) & access_T_CP_0_elements(243) & access_T_CP_0_elements(525);
      gj_access_T_cp_element_group_523 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(523), clk => clk, reset => reset); --
    end block;
    -- CP-element group 524:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: marked-predecessors 
    -- CP-element group 524: 	528 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	526 
    -- CP-element group 524:  members (3) 
      -- CP-element group 524: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_Update/req
      -- CP-element group 524: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_Update/$entry
      -- CP-element group 524: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_update_start_
      -- 
    req_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(524), ack => W_send1_4_752_delayed_14_0_788_inst_req_1); -- 
    access_T_cp_element_group_524: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_524"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(528);
      gj_access_T_cp_element_group_524 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(524), clk => clk, reset => reset); --
    end block;
    -- CP-element group 525:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	523 
    -- CP-element group 525: successors 
    -- CP-element group 525: marked-successors 
    -- CP-element group 525: 	313 
    -- CP-element group 525: 	77 
    -- CP-element group 525: 	523 
    -- CP-element group 525: 	239 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_Sample/ack
      -- CP-element group 525: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_Sample/$exit
      -- CP-element group 525: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_sample_completed_
      -- 
    ack_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send1_4_752_delayed_14_0_788_inst_ack_0, ack => access_T_CP_0_elements(525)); -- 
    -- CP-element group 526:  transition  input  bypass  pipeline-parent 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	524 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	527 
    -- CP-element group 526:  members (3) 
      -- CP-element group 526: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_Update/ack
      -- CP-element group 526: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_Update/$exit
      -- CP-element group 526: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_790_update_completed_
      -- 
    ack_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 526_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send1_4_752_delayed_14_0_788_inst_ack_1, ack => access_T_CP_0_elements(526)); -- 
    -- CP-element group 527:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	510 
    -- CP-element group 527: 	526 
    -- CP-element group 527: marked-predecessors 
    -- CP-element group 527: 	550 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	528 
    -- CP-element group 527:  members (3) 
      -- CP-element group 527: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_Sample/$entry
      -- CP-element group 527: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_Sample/req
      -- CP-element group 527: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_sample_start_
      -- 
    req_1774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(527), ack => WPIPE_input_pipe4_792_inst_req_0); -- 
    access_T_cp_element_group_527: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_527"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(510) & access_T_CP_0_elements(526) & access_T_CP_0_elements(550);
      gj_access_T_cp_element_group_527 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(527), clk => clk, reset => reset); --
    end block;
    -- CP-element group 528:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	527 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	529 
    -- CP-element group 528: marked-successors 
    -- CP-element group 528: 	508 
    -- CP-element group 528: 	524 
    -- CP-element group 528:  members (6) 
      -- CP-element group 528: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_Sample/ack
      -- CP-element group 528: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_Sample/$exit
      -- CP-element group 528: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_update_start_
      -- CP-element group 528: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_sample_completed_
      -- CP-element group 528: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_Update/req
      -- CP-element group 528: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_Update/$entry
      -- 
    ack_1775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_792_inst_ack_0, ack => access_T_CP_0_elements(528)); -- 
    req_1779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(528), ack => WPIPE_input_pipe4_792_inst_req_1); -- 
    -- CP-element group 529:  transition  input  bypass  pipeline-parent 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	528 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	534 
    -- CP-element group 529:  members (3) 
      -- CP-element group 529: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_update_completed_
      -- CP-element group 529: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_Update/ack
      -- CP-element group 529: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_792_Update/$exit
      -- 
    ack_1780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 529_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_792_inst_ack_1, ack => access_T_CP_0_elements(529)); -- 
    -- CP-element group 530:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	165 
    -- CP-element group 530: 	317 
    -- CP-element group 530: 	81 
    -- CP-element group 530: 	243 
    -- CP-element group 530: marked-predecessors 
    -- CP-element group 530: 	532 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	532 
    -- CP-element group 530:  members (3) 
      -- CP-element group 530: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_sample_start_
      -- CP-element group 530: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_Sample/$entry
      -- CP-element group 530: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_Sample/req
      -- 
    req_1788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(530), ack => W_send2_4_756_delayed_14_0_795_inst_req_0); -- 
    access_T_cp_element_group_530: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_530"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(165) & access_T_CP_0_elements(317) & access_T_CP_0_elements(81) & access_T_CP_0_elements(243) & access_T_CP_0_elements(532);
      gj_access_T_cp_element_group_530 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(530), clk => clk, reset => reset); --
    end block;
    -- CP-element group 531:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: marked-predecessors 
    -- CP-element group 531: 	535 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	533 
    -- CP-element group 531:  members (3) 
      -- CP-element group 531: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_Update/req
      -- CP-element group 531: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_Update/$entry
      -- CP-element group 531: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_update_start_
      -- 
    req_1793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(531), ack => W_send2_4_756_delayed_14_0_795_inst_req_1); -- 
    access_T_cp_element_group_531: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_531"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(535);
      gj_access_T_cp_element_group_531 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(531), clk => clk, reset => reset); --
    end block;
    -- CP-element group 532:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	530 
    -- CP-element group 532: successors 
    -- CP-element group 532: marked-successors 
    -- CP-element group 532: 	161 
    -- CP-element group 532: 	313 
    -- CP-element group 532: 	77 
    -- CP-element group 532: 	530 
    -- CP-element group 532: 	239 
    -- CP-element group 532:  members (3) 
      -- CP-element group 532: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_Sample/$exit
      -- CP-element group 532: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_Sample/ack
      -- CP-element group 532: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_sample_completed_
      -- 
    ack_1789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 532_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send2_4_756_delayed_14_0_795_inst_ack_0, ack => access_T_CP_0_elements(532)); -- 
    -- CP-element group 533:  transition  input  bypass  pipeline-parent 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	531 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	534 
    -- CP-element group 533:  members (3) 
      -- CP-element group 533: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_Update/$exit
      -- CP-element group 533: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_update_completed_
      -- CP-element group 533: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_797_Update/ack
      -- 
    ack_1794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 533_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send2_4_756_delayed_14_0_795_inst_ack_1, ack => access_T_CP_0_elements(533)); -- 
    -- CP-element group 534:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	514 
    -- CP-element group 534: 	529 
    -- CP-element group 534: 	533 
    -- CP-element group 534: marked-predecessors 
    -- CP-element group 534: 	536 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	535 
    -- CP-element group 534:  members (3) 
      -- CP-element group 534: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_sample_start_
      -- CP-element group 534: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_Sample/$entry
      -- CP-element group 534: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_Sample/req
      -- 
    req_1802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(534), ack => WPIPE_input_pipe4_799_inst_req_0); -- 
    access_T_cp_element_group_534: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_534"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(514) & access_T_CP_0_elements(529) & access_T_CP_0_elements(533) & access_T_CP_0_elements(536);
      gj_access_T_cp_element_group_534 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(534), clk => clk, reset => reset); --
    end block;
    -- CP-element group 535:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	534 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	536 
    -- CP-element group 535: marked-successors 
    -- CP-element group 535: 	512 
    -- CP-element group 535: 	531 
    -- CP-element group 535:  members (6) 
      -- CP-element group 535: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_sample_completed_
      -- CP-element group 535: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_update_start_
      -- CP-element group 535: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_Sample/$exit
      -- CP-element group 535: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_Sample/ack
      -- CP-element group 535: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_Update/$entry
      -- CP-element group 535: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_Update/req
      -- 
    ack_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 535_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_799_inst_ack_0, ack => access_T_CP_0_elements(535)); -- 
    req_1807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(535), ack => WPIPE_input_pipe4_799_inst_req_1); -- 
    -- CP-element group 536:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	535 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	541 
    -- CP-element group 536: marked-successors 
    -- CP-element group 536: 	534 
    -- CP-element group 536:  members (3) 
      -- CP-element group 536: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_update_completed_
      -- CP-element group 536: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_Update/$exit
      -- CP-element group 536: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_799_Update/ack
      -- 
    ack_1808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 536_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_799_inst_ack_1, ack => access_T_CP_0_elements(536)); -- 
    -- CP-element group 537:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	165 
    -- CP-element group 537: 	317 
    -- CP-element group 537: 	81 
    -- CP-element group 537: 	243 
    -- CP-element group 537: marked-predecessors 
    -- CP-element group 537: 	539 
    -- CP-element group 537: successors 
    -- CP-element group 537: 	539 
    -- CP-element group 537:  members (3) 
      -- CP-element group 537: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_sample_start_
      -- CP-element group 537: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_Sample/$entry
      -- CP-element group 537: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_Sample/req
      -- 
    req_1816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(537), ack => W_send3_4_760_delayed_14_0_802_inst_req_0); -- 
    access_T_cp_element_group_537: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_537"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(165) & access_T_CP_0_elements(317) & access_T_CP_0_elements(81) & access_T_CP_0_elements(243) & access_T_CP_0_elements(539);
      gj_access_T_cp_element_group_537 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(537), clk => clk, reset => reset); --
    end block;
    -- CP-element group 538:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: marked-predecessors 
    -- CP-element group 538: 	542 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	540 
    -- CP-element group 538:  members (3) 
      -- CP-element group 538: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_update_start_
      -- CP-element group 538: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_Update/$entry
      -- CP-element group 538: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_Update/req
      -- 
    req_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(538), ack => W_send3_4_760_delayed_14_0_802_inst_req_1); -- 
    access_T_cp_element_group_538: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_538"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(542);
      gj_access_T_cp_element_group_538 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(538), clk => clk, reset => reset); --
    end block;
    -- CP-element group 539:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	537 
    -- CP-element group 539: successors 
    -- CP-element group 539: marked-successors 
    -- CP-element group 539: 	161 
    -- CP-element group 539: 	313 
    -- CP-element group 539: 	77 
    -- CP-element group 539: 	537 
    -- CP-element group 539: 	239 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_sample_completed_
      -- CP-element group 539: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_Sample/$exit
      -- CP-element group 539: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_Sample/ack
      -- 
    ack_1817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 539_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send3_4_760_delayed_14_0_802_inst_ack_0, ack => access_T_CP_0_elements(539)); -- 
    -- CP-element group 540:  transition  input  bypass  pipeline-parent 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	538 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	541 
    -- CP-element group 540:  members (3) 
      -- CP-element group 540: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_update_completed_
      -- CP-element group 540: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_Update/$exit
      -- CP-element group 540: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_804_Update/ack
      -- 
    ack_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send3_4_760_delayed_14_0_802_inst_ack_1, ack => access_T_CP_0_elements(540)); -- 
    -- CP-element group 541:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	518 
    -- CP-element group 541: 	536 
    -- CP-element group 541: 	540 
    -- CP-element group 541: marked-predecessors 
    -- CP-element group 541: 	543 
    -- CP-element group 541: successors 
    -- CP-element group 541: 	542 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_sample_start_
      -- CP-element group 541: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_Sample/$entry
      -- CP-element group 541: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_Sample/req
      -- 
    req_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(541), ack => WPIPE_input_pipe4_806_inst_req_0); -- 
    access_T_cp_element_group_541: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_541"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(518) & access_T_CP_0_elements(536) & access_T_CP_0_elements(540) & access_T_CP_0_elements(543);
      gj_access_T_cp_element_group_541 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(541), clk => clk, reset => reset); --
    end block;
    -- CP-element group 542:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	541 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	543 
    -- CP-element group 542: marked-successors 
    -- CP-element group 542: 	516 
    -- CP-element group 542: 	538 
    -- CP-element group 542:  members (6) 
      -- CP-element group 542: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_sample_completed_
      -- CP-element group 542: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_update_start_
      -- CP-element group 542: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_Sample/$exit
      -- CP-element group 542: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_Sample/ack
      -- CP-element group 542: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_Update/$entry
      -- CP-element group 542: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_Update/req
      -- 
    ack_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 542_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_806_inst_ack_0, ack => access_T_CP_0_elements(542)); -- 
    req_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(542), ack => WPIPE_input_pipe4_806_inst_req_1); -- 
    -- CP-element group 543:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	542 
    -- CP-element group 543: successors 
    -- CP-element group 543: 	548 
    -- CP-element group 543: marked-successors 
    -- CP-element group 543: 	541 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_update_completed_
      -- CP-element group 543: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_Update/$exit
      -- CP-element group 543: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_806_Update/ack
      -- 
    ack_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 543_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_806_inst_ack_1, ack => access_T_CP_0_elements(543)); -- 
    -- CP-element group 544:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	165 
    -- CP-element group 544: 	317 
    -- CP-element group 544: 	243 
    -- CP-element group 544: marked-predecessors 
    -- CP-element group 544: 	546 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	546 
    -- CP-element group 544:  members (3) 
      -- CP-element group 544: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_sample_start_
      -- CP-element group 544: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_Sample/$entry
      -- CP-element group 544: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_Sample/req
      -- 
    req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(544), ack => W_send4_4_764_delayed_14_0_809_inst_req_0); -- 
    access_T_cp_element_group_544: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_544"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(165) & access_T_CP_0_elements(317) & access_T_CP_0_elements(243) & access_T_CP_0_elements(546);
      gj_access_T_cp_element_group_544 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(544), clk => clk, reset => reset); --
    end block;
    -- CP-element group 545:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: marked-predecessors 
    -- CP-element group 545: 	549 
    -- CP-element group 545: successors 
    -- CP-element group 545: 	547 
    -- CP-element group 545:  members (3) 
      -- CP-element group 545: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_update_start_
      -- CP-element group 545: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_Update/$entry
      -- CP-element group 545: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_Update/req
      -- 
    req_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(545), ack => W_send4_4_764_delayed_14_0_809_inst_req_1); -- 
    access_T_cp_element_group_545: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_545"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(549);
      gj_access_T_cp_element_group_545 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(545), clk => clk, reset => reset); --
    end block;
    -- CP-element group 546:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	544 
    -- CP-element group 546: successors 
    -- CP-element group 546: marked-successors 
    -- CP-element group 546: 	161 
    -- CP-element group 546: 	313 
    -- CP-element group 546: 	544 
    -- CP-element group 546: 	239 
    -- CP-element group 546:  members (3) 
      -- CP-element group 546: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_sample_completed_
      -- CP-element group 546: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_Sample/$exit
      -- CP-element group 546: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_Sample/ack
      -- 
    ack_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 546_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send4_4_764_delayed_14_0_809_inst_ack_0, ack => access_T_CP_0_elements(546)); -- 
    -- CP-element group 547:  transition  input  bypass  pipeline-parent 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	545 
    -- CP-element group 547: successors 
    -- CP-element group 547: 	548 
    -- CP-element group 547:  members (3) 
      -- CP-element group 547: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_update_completed_
      -- CP-element group 547: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_Update/$exit
      -- CP-element group 547: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_811_Update/ack
      -- 
    ack_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 547_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send4_4_764_delayed_14_0_809_inst_ack_1, ack => access_T_CP_0_elements(547)); -- 
    -- CP-element group 548:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	522 
    -- CP-element group 548: 	543 
    -- CP-element group 548: 	547 
    -- CP-element group 548: marked-predecessors 
    -- CP-element group 548: 	550 
    -- CP-element group 548: successors 
    -- CP-element group 548: 	549 
    -- CP-element group 548:  members (3) 
      -- CP-element group 548: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_sample_start_
      -- CP-element group 548: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_Sample/$entry
      -- CP-element group 548: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_Sample/req
      -- 
    req_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(548), ack => WPIPE_input_pipe4_813_inst_req_0); -- 
    access_T_cp_element_group_548: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_548"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(522) & access_T_CP_0_elements(543) & access_T_CP_0_elements(547) & access_T_CP_0_elements(550);
      gj_access_T_cp_element_group_548 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(548), clk => clk, reset => reset); --
    end block;
    -- CP-element group 549:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	548 
    -- CP-element group 549: successors 
    -- CP-element group 549: 	550 
    -- CP-element group 549: marked-successors 
    -- CP-element group 549: 	520 
    -- CP-element group 549: 	545 
    -- CP-element group 549:  members (6) 
      -- CP-element group 549: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_sample_completed_
      -- CP-element group 549: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_update_start_
      -- CP-element group 549: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_Sample/$exit
      -- CP-element group 549: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_Sample/ack
      -- CP-element group 549: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_Update/$entry
      -- CP-element group 549: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_Update/req
      -- 
    ack_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 549_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_813_inst_ack_0, ack => access_T_CP_0_elements(549)); -- 
    req_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(549), ack => WPIPE_input_pipe4_813_inst_req_1); -- 
    -- CP-element group 550:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	549 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	552 
    -- CP-element group 550: marked-successors 
    -- CP-element group 550: 	527 
    -- CP-element group 550: 	548 
    -- CP-element group 550:  members (3) 
      -- CP-element group 550: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_update_completed_
      -- CP-element group 550: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_Update/$exit
      -- CP-element group 550: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_813_Update/ack
      -- 
    ack_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 550_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_813_inst_ack_1, ack => access_T_CP_0_elements(550)); -- 
    -- CP-element group 551:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	9 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	10 
    -- CP-element group 551:  members (1) 
      -- CP-element group 551: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(551) is a control-delay.
    cp_element_551_delay: control_delay_element  generic map(name => " 551_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(551), clk => clk, reset =>reset);
    -- CP-element group 552:  join  transition  bypass  pipeline-parent 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	495 
    -- CP-element group 552: 	499 
    -- CP-element group 552: 	440 
    -- CP-element group 552: 	444 
    -- CP-element group 552: 	389 
    -- CP-element group 552: 	550 
    -- CP-element group 552: 	385 
    -- CP-element group 552: 	12 
    -- CP-element group 552: 	334 
    -- CP-element group 552: successors 
    -- CP-element group 552: 	6 
    -- CP-element group 552:  members (1) 
      -- CP-element group 552: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/$exit
      -- 
    access_T_cp_element_group_552: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_552"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= access_T_CP_0_elements(495) & access_T_CP_0_elements(499) & access_T_CP_0_elements(440) & access_T_CP_0_elements(444) & access_T_CP_0_elements(389) & access_T_CP_0_elements(550) & access_T_CP_0_elements(385) & access_T_CP_0_elements(12) & access_T_CP_0_elements(334);
      gj_access_T_cp_element_group_552 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(552), clk => clk, reset => reset); --
    end block;
    -- CP-element group 553:  transition  input  bypass  pipeline-parent 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	5 
    -- CP-element group 553: successors 
    -- CP-element group 553:  members (2) 
      -- CP-element group 553: 	 branch_block_stmt_29/do_while_stmt_42/loop_exit/$exit
      -- CP-element group 553: 	 branch_block_stmt_29/do_while_stmt_42/loop_exit/ack
      -- 
    ack_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_42_branch_ack_0, ack => access_T_CP_0_elements(553)); -- 
    -- CP-element group 554:  transition  input  bypass  pipeline-parent 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	5 
    -- CP-element group 554: successors 
    -- CP-element group 554:  members (2) 
      -- CP-element group 554: 	 branch_block_stmt_29/do_while_stmt_42/loop_taken/$exit
      -- CP-element group 554: 	 branch_block_stmt_29/do_while_stmt_42/loop_taken/ack
      -- 
    ack_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 554_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_42_branch_ack_1, ack => access_T_CP_0_elements(554)); -- 
    -- CP-element group 555:  transition  bypass  pipeline-parent 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	3 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	1 
    -- CP-element group 555:  members (1) 
      -- CP-element group 555: 	 branch_block_stmt_29/do_while_stmt_42/$exit
      -- 
    access_T_CP_0_elements(555) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_42_terminator_1874: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_42_terminator_1874", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(554),loop_terminate => access_T_CP_0_elements(553),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_44_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(23);
      access_T_CP_0_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(26);
      access_T_CP_0_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(32);
      access_T_CP_0_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(33);
      access_T_CP_0_elements(22) <= phi_mux_reqs(1);
      phi_stmt_44_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_44_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(17), 
          phi_sample_ack => access_T_CP_0_elements(18), 
          phi_update_req => access_T_CP_0_elements(19), 
          phi_update_ack => access_T_CP_0_elements(20), 
          phi_mux_ack => access_T_CP_0_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_49_phi_seq_132_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(48);
      access_T_CP_0_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(53);
      access_T_CP_0_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(54);
      access_T_CP_0_elements(43) <= phi_mux_reqs(1);
      phi_stmt_49_phi_seq_132 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_49_phi_seq_132") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(36), 
          phi_sample_ack => access_T_CP_0_elements(37), 
          phi_update_req => access_T_CP_0_elements(38), 
          phi_update_ack => access_T_CP_0_elements(39), 
          phi_mux_ack => access_T_CP_0_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_54_phi_seq_186_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(61);
      access_T_CP_0_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(68);
      access_T_CP_0_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(69);
      access_T_CP_0_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(63);
      access_T_CP_0_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(74);
      access_T_CP_0_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(75);
      access_T_CP_0_elements(64) <= phi_mux_reqs(1);
      phi_stmt_54_phi_seq_186 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_54_phi_seq_186") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(57), 
          phi_sample_ack => access_T_CP_0_elements(58), 
          phi_update_req => access_T_CP_0_elements(59), 
          phi_update_ack => access_T_CP_0_elements(60), 
          phi_mux_ack => access_T_CP_0_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_59_phi_seq_240_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(84);
      access_T_CP_0_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(91);
      access_T_CP_0_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(92);
      access_T_CP_0_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(82);
      access_T_CP_0_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(95);
      access_T_CP_0_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(96);
      access_T_CP_0_elements(83) <= phi_mux_reqs(1);
      phi_stmt_59_phi_seq_240 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_59_phi_seq_240") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(78), 
          phi_sample_ack => access_T_CP_0_elements(79), 
          phi_update_req => access_T_CP_0_elements(80), 
          phi_update_ack => access_T_CP_0_elements(81), 
          phi_mux_ack => access_T_CP_0_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_66_phi_seq_294_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(105);
      access_T_CP_0_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(112);
      access_T_CP_0_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(113);
      access_T_CP_0_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(103);
      access_T_CP_0_elements(114)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(115)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(117);
      access_T_CP_0_elements(104) <= phi_mux_reqs(1);
      phi_stmt_66_phi_seq_294 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_66_phi_seq_294") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(99), 
          phi_sample_ack => access_T_CP_0_elements(100), 
          phi_update_req => access_T_CP_0_elements(101), 
          phi_update_ack => access_T_CP_0_elements(102), 
          phi_mux_ack => access_T_CP_0_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_71_phi_seq_348_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(126);
      access_T_CP_0_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(133);
      access_T_CP_0_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(134);
      access_T_CP_0_elements(127) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(124);
      access_T_CP_0_elements(135)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(136)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(138);
      access_T_CP_0_elements(125) <= phi_mux_reqs(1);
      phi_stmt_71_phi_seq_348 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_71_phi_seq_348") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(120), 
          phi_sample_ack => access_T_CP_0_elements(121), 
          phi_update_req => access_T_CP_0_elements(122), 
          phi_update_ack => access_T_CP_0_elements(123), 
          phi_mux_ack => access_T_CP_0_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_76_phi_seq_402_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(147);
      access_T_CP_0_elements(150)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(154);
      access_T_CP_0_elements(151)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(155);
      access_T_CP_0_elements(148) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(145);
      access_T_CP_0_elements(156)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(158);
      access_T_CP_0_elements(157)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(159);
      access_T_CP_0_elements(146) <= phi_mux_reqs(1);
      phi_stmt_76_phi_seq_402 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_76_phi_seq_402") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(141), 
          phi_sample_ack => access_T_CP_0_elements(142), 
          phi_update_req => access_T_CP_0_elements(143), 
          phi_update_ack => access_T_CP_0_elements(144), 
          phi_mux_ack => access_T_CP_0_elements(149), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_81_phi_seq_456_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(168);
      access_T_CP_0_elements(171)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(175);
      access_T_CP_0_elements(172)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(176);
      access_T_CP_0_elements(169) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(166);
      access_T_CP_0_elements(177)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(179);
      access_T_CP_0_elements(178)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(180);
      access_T_CP_0_elements(167) <= phi_mux_reqs(1);
      phi_stmt_81_phi_seq_456 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_81_phi_seq_456") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(162), 
          phi_sample_ack => access_T_CP_0_elements(163), 
          phi_update_req => access_T_CP_0_elements(164), 
          phi_update_ack => access_T_CP_0_elements(165), 
          phi_mux_ack => access_T_CP_0_elements(170), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_86_phi_seq_500_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(187);
      access_T_CP_0_elements(192)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(194);
      access_T_CP_0_elements(193)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(195);
      access_T_CP_0_elements(188) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(189);
      access_T_CP_0_elements(196)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(196);
      access_T_CP_0_elements(197)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(198);
      access_T_CP_0_elements(190) <= phi_mux_reqs(1);
      phi_stmt_86_phi_seq_500 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_86_phi_seq_500") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(183), 
          phi_sample_ack => access_T_CP_0_elements(184), 
          phi_update_req => access_T_CP_0_elements(185), 
          phi_update_ack => access_T_CP_0_elements(186), 
          phi_mux_ack => access_T_CP_0_elements(191), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_91_phi_seq_544_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(208);
      access_T_CP_0_elements(211)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(211);
      access_T_CP_0_elements(212)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(213);
      access_T_CP_0_elements(209) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(206);
      access_T_CP_0_elements(215)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(217);
      access_T_CP_0_elements(216)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(218);
      access_T_CP_0_elements(207) <= phi_mux_reqs(1);
      phi_stmt_91_phi_seq_544 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_91_phi_seq_544") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(202), 
          phi_sample_ack => access_T_CP_0_elements(203), 
          phi_update_req => access_T_CP_0_elements(204), 
          phi_update_ack => access_T_CP_0_elements(205), 
          phi_mux_ack => access_T_CP_0_elements(210), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_96_phi_seq_588_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(227);
      access_T_CP_0_elements(230)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(230);
      access_T_CP_0_elements(231)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(232);
      access_T_CP_0_elements(228) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(225);
      access_T_CP_0_elements(234)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(236);
      access_T_CP_0_elements(235)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(237);
      access_T_CP_0_elements(226) <= phi_mux_reqs(1);
      phi_stmt_96_phi_seq_588 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_96_phi_seq_588") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(221), 
          phi_sample_ack => access_T_CP_0_elements(222), 
          phi_update_req => access_T_CP_0_elements(223), 
          phi_update_ack => access_T_CP_0_elements(224), 
          phi_mux_ack => access_T_CP_0_elements(229), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_101_phi_seq_632_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(246);
      access_T_CP_0_elements(249)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(249);
      access_T_CP_0_elements(250)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(251);
      access_T_CP_0_elements(247) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(244);
      access_T_CP_0_elements(253)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(255);
      access_T_CP_0_elements(254)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(256);
      access_T_CP_0_elements(245) <= phi_mux_reqs(1);
      phi_stmt_101_phi_seq_632 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_101_phi_seq_632") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(240), 
          phi_sample_ack => access_T_CP_0_elements(241), 
          phi_update_req => access_T_CP_0_elements(242), 
          phi_update_ack => access_T_CP_0_elements(243), 
          phi_mux_ack => access_T_CP_0_elements(248), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_106_phi_seq_676_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(265);
      access_T_CP_0_elements(268)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(268);
      access_T_CP_0_elements(269)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(270);
      access_T_CP_0_elements(266) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(263);
      access_T_CP_0_elements(272)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(274);
      access_T_CP_0_elements(273)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(275);
      access_T_CP_0_elements(264) <= phi_mux_reqs(1);
      phi_stmt_106_phi_seq_676 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_106_phi_seq_676") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(259), 
          phi_sample_ack => access_T_CP_0_elements(260), 
          phi_update_req => access_T_CP_0_elements(261), 
          phi_update_ack => access_T_CP_0_elements(262), 
          phi_mux_ack => access_T_CP_0_elements(267), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_111_phi_seq_720_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(282);
      access_T_CP_0_elements(285)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(285);
      access_T_CP_0_elements(286)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(287);
      access_T_CP_0_elements(283) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(280);
      access_T_CP_0_elements(289)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(291);
      access_T_CP_0_elements(290)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(292);
      access_T_CP_0_elements(281) <= phi_mux_reqs(1);
      phi_stmt_111_phi_seq_720 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_111_phi_seq_720") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(278), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(279), 
          phi_mux_ack => access_T_CP_0_elements(284), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_116_phi_seq_764_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(301);
      access_T_CP_0_elements(304)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(304);
      access_T_CP_0_elements(305)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(306);
      access_T_CP_0_elements(302) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(299);
      access_T_CP_0_elements(308)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(310);
      access_T_CP_0_elements(309)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(311);
      access_T_CP_0_elements(300) <= phi_mux_reqs(1);
      phi_stmt_116_phi_seq_764 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_116_phi_seq_764") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(295), 
          phi_sample_ack => access_T_CP_0_elements(296), 
          phi_update_req => access_T_CP_0_elements(297), 
          phi_update_ack => access_T_CP_0_elements(298), 
          phi_mux_ack => access_T_CP_0_elements(303), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_121_phi_seq_808_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(320);
      access_T_CP_0_elements(323)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(323);
      access_T_CP_0_elements(324)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(325);
      access_T_CP_0_elements(321) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(318);
      access_T_CP_0_elements(327)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(329);
      access_T_CP_0_elements(328)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(330);
      access_T_CP_0_elements(319) <= phi_mux_reqs(1);
      phi_stmt_121_phi_seq_808 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_121_phi_seq_808") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(314), 
          phi_sample_ack => access_T_CP_0_elements(315), 
          phi_update_req => access_T_CP_0_elements(316), 
          phi_update_ack => access_T_CP_0_elements(317), 
          phi_mux_ack => access_T_CP_0_elements(322), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_190_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_362_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_534_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_706_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_181_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_199_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_353_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_371_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_525_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_543_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_63_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_697_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_715_wire : std_logic_vector(31 downto 0);
    signal AND_u1_u1_237_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_243_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_253_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_259_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_409_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_415_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_425_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_431_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_581_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_587_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_597_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_603_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_753_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_759_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_769_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_775_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_225_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_397_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_569_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_741_wire : std_logic_vector(0 downto 0);
    signal LSHR_u64_u64_137_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_137_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_137_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_310_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_310_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_310_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_482_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_482_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_482_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_654_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_654_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_654_wire : std_logic_vector(63 downto 0);
    signal MUL_u16_u16_34_wire : std_logic_vector(15 downto 0);
    signal MUX_183_wire : std_logic_vector(31 downto 0);
    signal MUX_207_wire : std_logic_vector(63 downto 0);
    signal MUX_208_wire : std_logic_vector(63 downto 0);
    signal MUX_355_wire : std_logic_vector(31 downto 0);
    signal MUX_379_wire : std_logic_vector(63 downto 0);
    signal MUX_380_wire : std_logic_vector(63 downto 0);
    signal MUX_527_wire : std_logic_vector(31 downto 0);
    signal MUX_551_wire : std_logic_vector(63 downto 0);
    signal MUX_552_wire : std_logic_vector(63 downto 0);
    signal MUX_699_wire : std_logic_vector(31 downto 0);
    signal MUX_723_wire : std_logic_vector(63 downto 0);
    signal MUX_724_wire : std_logic_vector(63 downto 0);
    signal NOT_u1_u1_227_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_239_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_255_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_399_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_411_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_427_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_571_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_583_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_599_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_743_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_755_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_771_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_228_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_244_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_260_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_269_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_400_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_416_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_432_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_441_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_572_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_588_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_604_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_613_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_744_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_760_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_776_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_785_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_819_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_822_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_823_wire : std_logic_vector(0 downto 0);
    signal SUB_u64_u64_205_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_377_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_549_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_721_wire : std_logic_vector(63 downto 0);
    signal UGT_u32_u1_242_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_258_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_268_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_414_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_430_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_440_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_586_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_602_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_612_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_758_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_774_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_784_wire : std_logic_vector(0 downto 0);
    signal ULE_u2_u1_236_wire : std_logic_vector(0 downto 0);
    signal ULE_u2_u1_252_wire : std_logic_vector(0 downto 0);
    signal ULE_u2_u1_408_wire : std_logic_vector(0 downto 0);
    signal ULE_u2_u1_424_wire : std_logic_vector(0 downto 0);
    signal ULE_u2_u1_580_wire : std_logic_vector(0 downto 0);
    signal ULE_u2_u1_596_wire : std_logic_vector(0 downto 0);
    signal ULE_u2_u1_752_wire : std_logic_vector(0 downto 0);
    signal ULE_u2_u1_768_wire : std_logic_vector(0 downto 0);
    signal address1_44 : std_logic_vector(63 downto 0);
    signal address2_49 : std_logic_vector(63 downto 0);
    signal address3_54 : std_logic_vector(63 downto 0);
    signal address4_59 : std_logic_vector(63 downto 0);
    signal array_obj_ref_138_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_138_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_138_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_138_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_138_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_138_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_311_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_311_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_311_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_311_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_311_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_311_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_483_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_483_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_483_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_483_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_483_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_483_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_655_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_655_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_655_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_655_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_655_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_655_root_address : std_logic_vector(13 downto 0);
    signal continue_flag1_220 : std_logic_vector(0 downto 0);
    signal continue_flag2_392 : std_logic_vector(0 downto 0);
    signal continue_flag3_564 : std_logic_vector(0 downto 0);
    signal continue_flag4_736 : std_logic_vector(0 downto 0);
    signal fetch_addr1_140 : std_logic_vector(31 downto 0);
    signal fetch_addr2_313 : std_logic_vector(31 downto 0);
    signal fetch_addr3_485 : std_logic_vector(31 downto 0);
    signal fetch_addr4_657 : std_logic_vector(31 downto 0);
    signal fv1_144 : std_logic_vector(63 downto 0);
    signal fv2_317 : std_logic_vector(63 downto 0);
    signal fv3_489 : std_logic_vector(63 downto 0);
    signal fv4_661 : std_logic_vector(63 downto 0);
    signal konst_129_wire_constant : std_logic_vector(31 downto 0);
    signal konst_136_wire_constant : std_logic_vector(63 downto 0);
    signal konst_171_wire_constant : std_logic_vector(31 downto 0);
    signal konst_189_wire_constant : std_logic_vector(15 downto 0);
    signal konst_202_wire_constant : std_logic_vector(63 downto 0);
    signal konst_206_wire_constant : std_logic_vector(63 downto 0);
    signal konst_224_wire_constant : std_logic_vector(1 downto 0);
    signal konst_235_wire_constant : std_logic_vector(1 downto 0);
    signal konst_241_wire_constant : std_logic_vector(31 downto 0);
    signal konst_251_wire_constant : std_logic_vector(1 downto 0);
    signal konst_257_wire_constant : std_logic_vector(31 downto 0);
    signal konst_267_wire_constant : std_logic_vector(31 downto 0);
    signal konst_302_wire_constant : std_logic_vector(31 downto 0);
    signal konst_309_wire_constant : std_logic_vector(63 downto 0);
    signal konst_343_wire_constant : std_logic_vector(31 downto 0);
    signal konst_361_wire_constant : std_logic_vector(15 downto 0);
    signal konst_374_wire_constant : std_logic_vector(63 downto 0);
    signal konst_378_wire_constant : std_logic_vector(63 downto 0);
    signal konst_396_wire_constant : std_logic_vector(1 downto 0);
    signal konst_39_wire_constant : std_logic_vector(31 downto 0);
    signal konst_407_wire_constant : std_logic_vector(1 downto 0);
    signal konst_413_wire_constant : std_logic_vector(31 downto 0);
    signal konst_423_wire_constant : std_logic_vector(1 downto 0);
    signal konst_429_wire_constant : std_logic_vector(31 downto 0);
    signal konst_439_wire_constant : std_logic_vector(31 downto 0);
    signal konst_474_wire_constant : std_logic_vector(31 downto 0);
    signal konst_481_wire_constant : std_logic_vector(63 downto 0);
    signal konst_515_wire_constant : std_logic_vector(31 downto 0);
    signal konst_533_wire_constant : std_logic_vector(15 downto 0);
    signal konst_546_wire_constant : std_logic_vector(63 downto 0);
    signal konst_550_wire_constant : std_logic_vector(63 downto 0);
    signal konst_568_wire_constant : std_logic_vector(1 downto 0);
    signal konst_579_wire_constant : std_logic_vector(1 downto 0);
    signal konst_585_wire_constant : std_logic_vector(31 downto 0);
    signal konst_595_wire_constant : std_logic_vector(1 downto 0);
    signal konst_601_wire_constant : std_logic_vector(31 downto 0);
    signal konst_611_wire_constant : std_logic_vector(31 downto 0);
    signal konst_646_wire_constant : std_logic_vector(31 downto 0);
    signal konst_653_wire_constant : std_logic_vector(63 downto 0);
    signal konst_687_wire_constant : std_logic_vector(31 downto 0);
    signal konst_705_wire_constant : std_logic_vector(15 downto 0);
    signal konst_718_wire_constant : std_logic_vector(63 downto 0);
    signal konst_722_wire_constant : std_logic_vector(63 downto 0);
    signal konst_740_wire_constant : std_logic_vector(1 downto 0);
    signal konst_751_wire_constant : std_logic_vector(1 downto 0);
    signal konst_757_wire_constant : std_logic_vector(31 downto 0);
    signal konst_767_wire_constant : std_logic_vector(1 downto 0);
    signal konst_773_wire_constant : std_logic_vector(31 downto 0);
    signal konst_783_wire_constant : std_logic_vector(31 downto 0);
    signal last2_1_165 : std_logic_vector(1 downto 0);
    signal last2_2_337 : std_logic_vector(1 downto 0);
    signal last2_3_509 : std_logic_vector(1 downto 0);
    signal last2_4_681 : std_logic_vector(1 downto 0);
    signal m2_factor_41 : std_logic_vector(31 downto 0);
    signal m_factor_36 : std_logic_vector(31 downto 0);
    signal mycounter1_66 : std_logic_vector(31 downto 0);
    signal mycounter2_71 : std_logic_vector(31 downto 0);
    signal mycounter3_76 : std_logic_vector(31 downto 0);
    signal mycounter4_81 : std_logic_vector(31 downto 0);
    signal n_address1_210 : std_logic_vector(63 downto 0);
    signal n_address1_210_48_buffered : std_logic_vector(63 downto 0);
    signal n_address2_382 : std_logic_vector(63 downto 0);
    signal n_address2_382_51_buffered : std_logic_vector(63 downto 0);
    signal n_address3_554 : std_logic_vector(63 downto 0);
    signal n_address3_554_56_buffered : std_logic_vector(63 downto 0);
    signal n_address4_726 : std_logic_vector(63 downto 0);
    signal n_address4_726_65_buffered : std_logic_vector(63 downto 0);
    signal n_mycounter1_185 : std_logic_vector(31 downto 0);
    signal n_mycounter1_185_70_buffered : std_logic_vector(31 downto 0);
    signal n_mycounter2_357 : std_logic_vector(31 downto 0);
    signal n_mycounter2_357_75_buffered : std_logic_vector(31 downto 0);
    signal n_mycounter3_529 : std_logic_vector(31 downto 0);
    signal n_mycounter3_529_80_buffered : std_logic_vector(31 downto 0);
    signal n_mycounter4_701 : std_logic_vector(31 downto 0);
    signal n_mycounter4_701_85_buffered : std_logic_vector(31 downto 0);
    signal n_row1_193 : std_logic_vector(15 downto 0);
    signal n_row1_193_88_buffered : std_logic_vector(15 downto 0);
    signal n_row2_365 : std_logic_vector(15 downto 0);
    signal n_row2_365_95_buffered : std_logic_vector(15 downto 0);
    signal n_row3_537 : std_logic_vector(15 downto 0);
    signal n_row3_537_100_buffered : std_logic_vector(15 downto 0);
    signal n_row4_709 : std_logic_vector(15 downto 0);
    signal n_row4_709_105_buffered : std_logic_vector(15 downto 0);
    signal n_start1_168 : std_logic_vector(0 downto 0);
    signal n_start1_168_110_buffered : std_logic_vector(0 downto 0);
    signal n_start2_340 : std_logic_vector(0 downto 0);
    signal n_start2_340_115_buffered : std_logic_vector(0 downto 0);
    signal n_start3_512 : std_logic_vector(0 downto 0);
    signal n_start3_512_120_buffered : std_logic_vector(0 downto 0);
    signal n_start4_684 : std_logic_vector(0 downto 0);
    signal n_start4_684_125_buffered : std_logic_vector(0 downto 0);
    signal next_row1_131 : std_logic_vector(0 downto 0);
    signal next_row2_304 : std_logic_vector(0 downto 0);
    signal next_row3_476 : std_logic_vector(0 downto 0);
    signal next_row4_648 : std_logic_vector(0 downto 0);
    signal ptr_deref_143_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_143_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_143_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_143_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_143_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_316_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_316_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_316_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_316_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_316_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_488_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_488_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_488_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_488_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_488_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_660_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_660_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_660_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_660_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_660_word_offset_0 : std_logic_vector(13 downto 0);
    signal row1_86 : std_logic_vector(15 downto 0);
    signal row2_91 : std_logic_vector(15 downto 0);
    signal row3_96 : std_logic_vector(15 downto 0);
    signal row4_101 : std_logic_vector(15 downto 0);
    signal send1_1_230 : std_logic_vector(0 downto 0);
    signal send1_1_272_delayed_14_0_274 : std_logic_vector(0 downto 0);
    signal send1_2_402 : std_logic_vector(0 downto 0);
    signal send1_2_432_delayed_14_0_446 : std_logic_vector(0 downto 0);
    signal send1_3_574 : std_logic_vector(0 downto 0);
    signal send1_3_592_delayed_14_0_618 : std_logic_vector(0 downto 0);
    signal send1_4_746 : std_logic_vector(0 downto 0);
    signal send1_4_752_delayed_14_0_790 : std_logic_vector(0 downto 0);
    signal send2_1_246 : std_logic_vector(0 downto 0);
    signal send2_1_276_delayed_14_0_281 : std_logic_vector(0 downto 0);
    signal send2_2_418 : std_logic_vector(0 downto 0);
    signal send2_2_436_delayed_14_0_453 : std_logic_vector(0 downto 0);
    signal send2_3_590 : std_logic_vector(0 downto 0);
    signal send2_3_596_delayed_14_0_625 : std_logic_vector(0 downto 0);
    signal send2_4_756_delayed_14_0_797 : std_logic_vector(0 downto 0);
    signal send2_4_762 : std_logic_vector(0 downto 0);
    signal send3_1_262 : std_logic_vector(0 downto 0);
    signal send3_1_280_delayed_14_0_288 : std_logic_vector(0 downto 0);
    signal send3_2_434 : std_logic_vector(0 downto 0);
    signal send3_2_440_delayed_14_0_460 : std_logic_vector(0 downto 0);
    signal send3_3_600_delayed_14_0_632 : std_logic_vector(0 downto 0);
    signal send3_3_606 : std_logic_vector(0 downto 0);
    signal send3_4_760_delayed_14_0_804 : std_logic_vector(0 downto 0);
    signal send3_4_778 : std_logic_vector(0 downto 0);
    signal send4_1_271 : std_logic_vector(0 downto 0);
    signal send4_1_284_delayed_14_0_295 : std_logic_vector(0 downto 0);
    signal send4_2_443 : std_logic_vector(0 downto 0);
    signal send4_2_444_delayed_14_0_467 : std_logic_vector(0 downto 0);
    signal send4_3_604_delayed_14_0_639 : std_logic_vector(0 downto 0);
    signal send4_3_615 : std_logic_vector(0 downto 0);
    signal send4_4_764_delayed_14_0_811 : std_logic_vector(0 downto 0);
    signal send4_4_787 : std_logic_vector(0 downto 0);
    signal send_flag1_215 : std_logic_vector(0 downto 0);
    signal send_flag2_387 : std_logic_vector(0 downto 0);
    signal send_flag3_559 : std_logic_vector(0 downto 0);
    signal send_flag4_731 : std_logic_vector(0 downto 0);
    signal start1_106 : std_logic_vector(0 downto 0);
    signal start2_111 : std_logic_vector(0 downto 0);
    signal start3_116 : std_logic_vector(0 downto 0);
    signal start4_121 : std_logic_vector(0 downto 0);
    signal tmp_cnt1_173 : std_logic_vector(31 downto 0);
    signal tmp_cnt2_345 : std_logic_vector(31 downto 0);
    signal tmp_cnt3_517 : std_logic_vector(31 downto 0);
    signal tmp_cnt4_689 : std_logic_vector(31 downto 0);
    signal type_cast_104_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_109_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_114_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_119_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_124_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_180_wire : std_logic_vector(31 downto 0);
    signal type_cast_200_wire : std_logic_vector(63 downto 0);
    signal type_cast_204_wire : std_logic_vector(63 downto 0);
    signal type_cast_352_wire : std_logic_vector(31 downto 0);
    signal type_cast_372_wire : std_logic_vector(63 downto 0);
    signal type_cast_376_wire : std_logic_vector(63 downto 0);
    signal type_cast_47_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_524_wire : std_logic_vector(31 downto 0);
    signal type_cast_53_wire : std_logic_vector(63 downto 0);
    signal type_cast_544_wire : std_logic_vector(63 downto 0);
    signal type_cast_548_wire : std_logic_vector(63 downto 0);
    signal type_cast_58_wire : std_logic_vector(63 downto 0);
    signal type_cast_64_wire : std_logic_vector(63 downto 0);
    signal type_cast_696_wire : std_logic_vector(31 downto 0);
    signal type_cast_69_wire : std_logic_vector(31 downto 0);
    signal type_cast_716_wire : std_logic_vector(63 downto 0);
    signal type_cast_720_wire : std_logic_vector(63 downto 0);
    signal type_cast_74_wire : std_logic_vector(31 downto 0);
    signal type_cast_79_wire : std_logic_vector(31 downto 0);
    signal type_cast_84_wire : std_logic_vector(31 downto 0);
    signal type_cast_90_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_99_wire_constant : std_logic_vector(15 downto 0);
    signal w_11_148 : std_logic_vector(15 downto 0);
    signal w_12_321 : std_logic_vector(15 downto 0);
    signal w_13_493 : std_logic_vector(15 downto 0);
    signal w_14_665 : std_logic_vector(15 downto 0);
    signal w_21_152 : std_logic_vector(15 downto 0);
    signal w_22_325 : std_logic_vector(15 downto 0);
    signal w_23_497 : std_logic_vector(15 downto 0);
    signal w_24_669 : std_logic_vector(15 downto 0);
    signal w_31_156 : std_logic_vector(15 downto 0);
    signal w_32_329 : std_logic_vector(15 downto 0);
    signal w_33_501 : std_logic_vector(15 downto 0);
    signal w_34_673 : std_logic_vector(15 downto 0);
    signal w_41_160 : std_logic_vector(15 downto 0);
    signal w_42_333 : std_logic_vector(15 downto 0);
    signal w_43_505 : std_logic_vector(15 downto 0);
    signal w_44_677 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_138_constant_part_of_offset <= "00000000000000";
    array_obj_ref_138_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_138_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_138_resized_base_address <= "00000000000000";
    array_obj_ref_311_constant_part_of_offset <= "00000000000000";
    array_obj_ref_311_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_311_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_311_resized_base_address <= "00000000000000";
    array_obj_ref_483_constant_part_of_offset <= "00000000000000";
    array_obj_ref_483_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_483_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_483_resized_base_address <= "00000000000000";
    array_obj_ref_655_constant_part_of_offset <= "00000000000000";
    array_obj_ref_655_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_655_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_655_resized_base_address <= "00000000000000";
    konst_129_wire_constant <= "00000000000000000000000000000100";
    konst_136_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_171_wire_constant <= "00000000000000000000000000000100";
    konst_189_wire_constant <= "0000000000000010";
    konst_202_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_206_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_224_wire_constant <= "00";
    konst_235_wire_constant <= "01";
    konst_241_wire_constant <= "00000000000000000000000000000001";
    konst_251_wire_constant <= "10";
    konst_257_wire_constant <= "00000000000000000000000000000010";
    konst_267_wire_constant <= "00000000000000000000000000000011";
    konst_302_wire_constant <= "00000000000000000000000000000100";
    konst_309_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_343_wire_constant <= "00000000000000000000000000000100";
    konst_361_wire_constant <= "0000000000000010";
    konst_374_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_378_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_396_wire_constant <= "00";
    konst_39_wire_constant <= "00000000000000000000000000000001";
    konst_407_wire_constant <= "01";
    konst_413_wire_constant <= "00000000000000000000000000000001";
    konst_423_wire_constant <= "10";
    konst_429_wire_constant <= "00000000000000000000000000000010";
    konst_439_wire_constant <= "00000000000000000000000000000011";
    konst_474_wire_constant <= "00000000000000000000000000000100";
    konst_481_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_515_wire_constant <= "00000000000000000000000000000100";
    konst_533_wire_constant <= "0000000000000010";
    konst_546_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_550_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_568_wire_constant <= "00";
    konst_579_wire_constant <= "01";
    konst_585_wire_constant <= "00000000000000000000000000000001";
    konst_595_wire_constant <= "10";
    konst_601_wire_constant <= "00000000000000000000000000000010";
    konst_611_wire_constant <= "00000000000000000000000000000011";
    konst_646_wire_constant <= "00000000000000000000000000000100";
    konst_653_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_687_wire_constant <= "00000000000000000000000000000100";
    konst_705_wire_constant <= "0000000000000010";
    konst_718_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_722_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_740_wire_constant <= "00";
    konst_751_wire_constant <= "01";
    konst_757_wire_constant <= "00000000000000000000000000000001";
    konst_767_wire_constant <= "10";
    konst_773_wire_constant <= "00000000000000000000000000000010";
    konst_783_wire_constant <= "00000000000000000000000000000011";
    ptr_deref_143_word_offset_0 <= "00000000000000";
    ptr_deref_316_word_offset_0 <= "00000000000000";
    ptr_deref_488_word_offset_0 <= "00000000000000";
    ptr_deref_660_word_offset_0 <= "00000000000000";
    type_cast_104_wire_constant <= "0000000000000001";
    type_cast_109_wire_constant <= "1";
    type_cast_114_wire_constant <= "1";
    type_cast_119_wire_constant <= "1";
    type_cast_124_wire_constant <= "1";
    type_cast_47_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_90_wire_constant <= "0000000000000000";
    type_cast_94_wire_constant <= "0000000000000000";
    type_cast_99_wire_constant <= "0000000000000000";
    phi_stmt_101: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_104_wire_constant & n_row4_709_105_buffered;
      req <= phi_stmt_101_req_0 & phi_stmt_101_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_101",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_101_ack_0,
          idata => idata,
          odata => row4_101,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_101
    phi_stmt_106: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_109_wire_constant & n_start1_168_110_buffered;
      req <= phi_stmt_106_req_0 & phi_stmt_106_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_106",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_106_ack_0,
          idata => idata,
          odata => start1_106,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_106
    phi_stmt_111: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_114_wire_constant & n_start2_340_115_buffered;
      req <= phi_stmt_111_req_0 & phi_stmt_111_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_111",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_111_ack_0,
          idata => idata,
          odata => start2_111,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_111
    phi_stmt_116: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_119_wire_constant & n_start3_512_120_buffered;
      req <= phi_stmt_116_req_0 & phi_stmt_116_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_116",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_116_ack_0,
          idata => idata,
          odata => start3_116,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_116
    phi_stmt_121: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_124_wire_constant & n_start4_684_125_buffered;
      req <= phi_stmt_121_req_0 & phi_stmt_121_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_121",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_121_ack_0,
          idata => idata,
          odata => start4_121,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_121
    phi_stmt_44: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_47_wire_constant & n_address1_210_48_buffered;
      req <= phi_stmt_44_req_0 & phi_stmt_44_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_44",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_44_ack_0,
          idata => idata,
          odata => address1_44,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_44
    phi_stmt_49: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address2_382_51_buffered & type_cast_53_wire;
      req <= phi_stmt_49_req_0 & phi_stmt_49_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_49",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_49_ack_0,
          idata => idata,
          odata => address2_49,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_49
    phi_stmt_54: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address3_554_56_buffered & type_cast_58_wire;
      req <= phi_stmt_54_req_0 & phi_stmt_54_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_54",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_54_ack_0,
          idata => idata,
          odata => address3_54,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_54
    phi_stmt_59: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_64_wire & n_address4_726_65_buffered;
      req <= phi_stmt_59_req_0 & phi_stmt_59_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_59",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_59_ack_0,
          idata => idata,
          odata => address4_59,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_59
    phi_stmt_66: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_69_wire & n_mycounter1_185_70_buffered;
      req <= phi_stmt_66_req_0 & phi_stmt_66_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_66",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_66_ack_0,
          idata => idata,
          odata => mycounter1_66,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_66
    phi_stmt_71: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_74_wire & n_mycounter2_357_75_buffered;
      req <= phi_stmt_71_req_0 & phi_stmt_71_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_71",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_71_ack_0,
          idata => idata,
          odata => mycounter2_71,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_71
    phi_stmt_76: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_79_wire & n_mycounter3_529_80_buffered;
      req <= phi_stmt_76_req_0 & phi_stmt_76_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_76",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_76_ack_0,
          idata => idata,
          odata => mycounter3_76,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_76
    phi_stmt_81: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_84_wire & n_mycounter4_701_85_buffered;
      req <= phi_stmt_81_req_0 & phi_stmt_81_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_81",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_81_ack_0,
          idata => idata,
          odata => mycounter4_81,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_81
    phi_stmt_86: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_row1_193_88_buffered & type_cast_90_wire_constant;
      req <= phi_stmt_86_req_0 & phi_stmt_86_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_86",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_86_ack_0,
          idata => idata,
          odata => row1_86,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_86
    phi_stmt_91: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_94_wire_constant & n_row2_365_95_buffered;
      req <= phi_stmt_91_req_0 & phi_stmt_91_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_91",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_91_ack_0,
          idata => idata,
          odata => row2_91,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_91
    phi_stmt_96: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_99_wire_constant & n_row3_537_100_buffered;
      req <= phi_stmt_96_req_0 & phi_stmt_96_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_96",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_96_ack_0,
          idata => idata,
          odata => row3_96,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_96
    -- flow-through select operator MUX_183_inst
    MUX_183_wire <= ADD_u32_u32_181_wire when (start1_106(0) /=  '0') else tmp_cnt1_173;
    -- flow-through select operator MUX_184_inst
    n_mycounter1_185 <= m_factor_36 when (next_row1_131(0) /=  '0') else MUX_183_wire;
    -- flow-through select operator MUX_192_inst
    n_row1_193 <= ADD_u16_u16_190_wire when (next_row1_131(0) /=  '0') else row1_86;
    -- flow-through select operator MUX_207_inst
    MUX_207_wire <= SUB_u64_u64_205_wire when (start1_106(0) /=  '0') else konst_206_wire_constant;
    -- flow-through select operator MUX_208_inst
    MUX_208_wire <= type_cast_200_wire when (next_row1_131(0) /=  '0') else MUX_207_wire;
    -- flow-through select operator MUX_355_inst
    MUX_355_wire <= ADD_u32_u32_353_wire when (start2_111(0) /=  '0') else tmp_cnt2_345;
    -- flow-through select operator MUX_356_inst
    n_mycounter2_357 <= m_factor_36 when (next_row2_304(0) /=  '0') else MUX_355_wire;
    -- flow-through select operator MUX_364_inst
    n_row2_365 <= ADD_u16_u16_362_wire when (next_row2_304(0) /=  '0') else row2_91;
    -- flow-through select operator MUX_379_inst
    MUX_379_wire <= SUB_u64_u64_377_wire when (start2_111(0) /=  '0') else konst_378_wire_constant;
    -- flow-through select operator MUX_380_inst
    MUX_380_wire <= type_cast_372_wire when (next_row2_304(0) /=  '0') else MUX_379_wire;
    -- flow-through select operator MUX_527_inst
    MUX_527_wire <= ADD_u32_u32_525_wire when (start3_116(0) /=  '0') else tmp_cnt3_517;
    -- flow-through select operator MUX_528_inst
    n_mycounter3_529 <= m_factor_36 when (next_row3_476(0) /=  '0') else MUX_527_wire;
    -- flow-through select operator MUX_536_inst
    n_row3_537 <= ADD_u16_u16_534_wire when (next_row3_476(0) /=  '0') else row3_96;
    -- flow-through select operator MUX_551_inst
    MUX_551_wire <= SUB_u64_u64_549_wire when (start3_116(0) /=  '0') else konst_550_wire_constant;
    -- flow-through select operator MUX_552_inst
    MUX_552_wire <= type_cast_544_wire when (next_row3_476(0) /=  '0') else MUX_551_wire;
    -- flow-through select operator MUX_699_inst
    MUX_699_wire <= ADD_u32_u32_697_wire when (start4_121(0) /=  '0') else tmp_cnt4_689;
    -- flow-through select operator MUX_700_inst
    n_mycounter4_701 <= m_factor_36 when (next_row4_648(0) /=  '0') else MUX_699_wire;
    -- flow-through select operator MUX_708_inst
    n_row4_709 <= ADD_u16_u16_706_wire when (next_row4_648(0) /=  '0') else row4_101;
    -- flow-through select operator MUX_723_inst
    MUX_723_wire <= SUB_u64_u64_721_wire when (start4_121(0) /=  '0') else konst_722_wire_constant;
    -- flow-through select operator MUX_724_inst
    MUX_724_wire <= type_cast_716_wire when (next_row4_648(0) /=  '0') else MUX_723_wire;
    slice_147_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_147_inst_req_0;
      slice_147_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_147_inst_req_1;
      slice_147_inst_ack_1<= update_ack(0);
      slice_147_inst: SliceSplitProtocol generic map(name => "slice_147_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv1_144, dout => w_11_148, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_151_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_151_inst_req_0;
      slice_151_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_151_inst_req_1;
      slice_151_inst_ack_1<= update_ack(0);
      slice_151_inst: SliceSplitProtocol generic map(name => "slice_151_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv1_144, dout => w_21_152, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_155_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_155_inst_req_0;
      slice_155_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_155_inst_req_1;
      slice_155_inst_ack_1<= update_ack(0);
      slice_155_inst: SliceSplitProtocol generic map(name => "slice_155_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv1_144, dout => w_31_156, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_159_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_159_inst_req_0;
      slice_159_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_159_inst_req_1;
      slice_159_inst_ack_1<= update_ack(0);
      slice_159_inst: SliceSplitProtocol generic map(name => "slice_159_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv1_144, dout => w_41_160, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_320_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_320_inst_req_0;
      slice_320_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_320_inst_req_1;
      slice_320_inst_ack_1<= update_ack(0);
      slice_320_inst: SliceSplitProtocol generic map(name => "slice_320_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv2_317, dout => w_12_321, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_324_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_324_inst_req_0;
      slice_324_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_324_inst_req_1;
      slice_324_inst_ack_1<= update_ack(0);
      slice_324_inst: SliceSplitProtocol generic map(name => "slice_324_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv2_317, dout => w_22_325, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_328_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_328_inst_req_0;
      slice_328_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_328_inst_req_1;
      slice_328_inst_ack_1<= update_ack(0);
      slice_328_inst: SliceSplitProtocol generic map(name => "slice_328_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv2_317, dout => w_32_329, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_332_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_332_inst_req_0;
      slice_332_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_332_inst_req_1;
      slice_332_inst_ack_1<= update_ack(0);
      slice_332_inst: SliceSplitProtocol generic map(name => "slice_332_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv2_317, dout => w_42_333, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_492_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_492_inst_req_0;
      slice_492_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_492_inst_req_1;
      slice_492_inst_ack_1<= update_ack(0);
      slice_492_inst: SliceSplitProtocol generic map(name => "slice_492_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv3_489, dout => w_13_493, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_496_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_496_inst_req_0;
      slice_496_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_496_inst_req_1;
      slice_496_inst_ack_1<= update_ack(0);
      slice_496_inst: SliceSplitProtocol generic map(name => "slice_496_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv3_489, dout => w_23_497, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_500_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_500_inst_req_0;
      slice_500_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_500_inst_req_1;
      slice_500_inst_ack_1<= update_ack(0);
      slice_500_inst: SliceSplitProtocol generic map(name => "slice_500_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv3_489, dout => w_33_501, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_504_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_504_inst_req_0;
      slice_504_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_504_inst_req_1;
      slice_504_inst_ack_1<= update_ack(0);
      slice_504_inst: SliceSplitProtocol generic map(name => "slice_504_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv3_489, dout => w_43_505, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_664_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_664_inst_req_0;
      slice_664_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_664_inst_req_1;
      slice_664_inst_ack_1<= update_ack(0);
      slice_664_inst: SliceSplitProtocol generic map(name => "slice_664_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv4_661, dout => w_14_665, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_668_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_668_inst_req_0;
      slice_668_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_668_inst_req_1;
      slice_668_inst_ack_1<= update_ack(0);
      slice_668_inst: SliceSplitProtocol generic map(name => "slice_668_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv4_661, dout => w_24_669, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_672_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_672_inst_req_0;
      slice_672_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_672_inst_req_1;
      slice_672_inst_ack_1<= update_ack(0);
      slice_672_inst: SliceSplitProtocol generic map(name => "slice_672_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv4_661, dout => w_34_673, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_676_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_676_inst_req_0;
      slice_676_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_676_inst_req_1;
      slice_676_inst_ack_1<= update_ack(0);
      slice_676_inst: SliceSplitProtocol generic map(name => "slice_676_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fv4_661, dout => w_44_677, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- interlock W_n_start1_166_inst
    process(next_row1_131) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := next_row1_131(0 downto 0);
      n_start1_168 <= tmp_var; -- 
    end process;
    -- interlock W_n_start2_338_inst
    process(next_row2_304) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := next_row2_304(0 downto 0);
      n_start2_340 <= tmp_var; -- 
    end process;
    -- interlock W_n_start3_510_inst
    process(next_row3_476) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := next_row3_476(0 downto 0);
      n_start3_512 <= tmp_var; -- 
    end process;
    -- interlock W_n_start4_682_inst
    process(next_row4_648) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := next_row4_648(0 downto 0);
      n_start4_684 <= tmp_var; -- 
    end process;
    W_send1_1_272_delayed_14_0_272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send1_1_272_delayed_14_0_272_inst_req_0;
      W_send1_1_272_delayed_14_0_272_inst_ack_0<= wack(0);
      rreq(0) <= W_send1_1_272_delayed_14_0_272_inst_req_1;
      W_send1_1_272_delayed_14_0_272_inst_ack_1<= rack(0);
      W_send1_1_272_delayed_14_0_272_inst : InterlockBuffer generic map ( -- 
        name => "W_send1_1_272_delayed_14_0_272_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send1_1_230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send1_1_272_delayed_14_0_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send1_2_432_delayed_14_0_444_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send1_2_432_delayed_14_0_444_inst_req_0;
      W_send1_2_432_delayed_14_0_444_inst_ack_0<= wack(0);
      rreq(0) <= W_send1_2_432_delayed_14_0_444_inst_req_1;
      W_send1_2_432_delayed_14_0_444_inst_ack_1<= rack(0);
      W_send1_2_432_delayed_14_0_444_inst : InterlockBuffer generic map ( -- 
        name => "W_send1_2_432_delayed_14_0_444_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send1_2_402,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send1_2_432_delayed_14_0_446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send1_3_592_delayed_14_0_616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send1_3_592_delayed_14_0_616_inst_req_0;
      W_send1_3_592_delayed_14_0_616_inst_ack_0<= wack(0);
      rreq(0) <= W_send1_3_592_delayed_14_0_616_inst_req_1;
      W_send1_3_592_delayed_14_0_616_inst_ack_1<= rack(0);
      W_send1_3_592_delayed_14_0_616_inst : InterlockBuffer generic map ( -- 
        name => "W_send1_3_592_delayed_14_0_616_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send1_3_574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send1_3_592_delayed_14_0_618,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send1_4_752_delayed_14_0_788_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send1_4_752_delayed_14_0_788_inst_req_0;
      W_send1_4_752_delayed_14_0_788_inst_ack_0<= wack(0);
      rreq(0) <= W_send1_4_752_delayed_14_0_788_inst_req_1;
      W_send1_4_752_delayed_14_0_788_inst_ack_1<= rack(0);
      W_send1_4_752_delayed_14_0_788_inst : InterlockBuffer generic map ( -- 
        name => "W_send1_4_752_delayed_14_0_788_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send1_4_746,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send1_4_752_delayed_14_0_790,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send2_1_276_delayed_14_0_279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send2_1_276_delayed_14_0_279_inst_req_0;
      W_send2_1_276_delayed_14_0_279_inst_ack_0<= wack(0);
      rreq(0) <= W_send2_1_276_delayed_14_0_279_inst_req_1;
      W_send2_1_276_delayed_14_0_279_inst_ack_1<= rack(0);
      W_send2_1_276_delayed_14_0_279_inst : InterlockBuffer generic map ( -- 
        name => "W_send2_1_276_delayed_14_0_279_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send2_1_246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send2_1_276_delayed_14_0_281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send2_2_436_delayed_14_0_451_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send2_2_436_delayed_14_0_451_inst_req_0;
      W_send2_2_436_delayed_14_0_451_inst_ack_0<= wack(0);
      rreq(0) <= W_send2_2_436_delayed_14_0_451_inst_req_1;
      W_send2_2_436_delayed_14_0_451_inst_ack_1<= rack(0);
      W_send2_2_436_delayed_14_0_451_inst : InterlockBuffer generic map ( -- 
        name => "W_send2_2_436_delayed_14_0_451_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send2_2_418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send2_2_436_delayed_14_0_453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send2_3_596_delayed_14_0_623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send2_3_596_delayed_14_0_623_inst_req_0;
      W_send2_3_596_delayed_14_0_623_inst_ack_0<= wack(0);
      rreq(0) <= W_send2_3_596_delayed_14_0_623_inst_req_1;
      W_send2_3_596_delayed_14_0_623_inst_ack_1<= rack(0);
      W_send2_3_596_delayed_14_0_623_inst : InterlockBuffer generic map ( -- 
        name => "W_send2_3_596_delayed_14_0_623_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send2_3_590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send2_3_596_delayed_14_0_625,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send2_4_756_delayed_14_0_795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send2_4_756_delayed_14_0_795_inst_req_0;
      W_send2_4_756_delayed_14_0_795_inst_ack_0<= wack(0);
      rreq(0) <= W_send2_4_756_delayed_14_0_795_inst_req_1;
      W_send2_4_756_delayed_14_0_795_inst_ack_1<= rack(0);
      W_send2_4_756_delayed_14_0_795_inst : InterlockBuffer generic map ( -- 
        name => "W_send2_4_756_delayed_14_0_795_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send2_4_762,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send2_4_756_delayed_14_0_797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send3_1_280_delayed_14_0_286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send3_1_280_delayed_14_0_286_inst_req_0;
      W_send3_1_280_delayed_14_0_286_inst_ack_0<= wack(0);
      rreq(0) <= W_send3_1_280_delayed_14_0_286_inst_req_1;
      W_send3_1_280_delayed_14_0_286_inst_ack_1<= rack(0);
      W_send3_1_280_delayed_14_0_286_inst : InterlockBuffer generic map ( -- 
        name => "W_send3_1_280_delayed_14_0_286_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send3_1_262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send3_1_280_delayed_14_0_288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send3_2_440_delayed_14_0_458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send3_2_440_delayed_14_0_458_inst_req_0;
      W_send3_2_440_delayed_14_0_458_inst_ack_0<= wack(0);
      rreq(0) <= W_send3_2_440_delayed_14_0_458_inst_req_1;
      W_send3_2_440_delayed_14_0_458_inst_ack_1<= rack(0);
      W_send3_2_440_delayed_14_0_458_inst : InterlockBuffer generic map ( -- 
        name => "W_send3_2_440_delayed_14_0_458_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send3_2_434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send3_2_440_delayed_14_0_460,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send3_3_600_delayed_14_0_630_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send3_3_600_delayed_14_0_630_inst_req_0;
      W_send3_3_600_delayed_14_0_630_inst_ack_0<= wack(0);
      rreq(0) <= W_send3_3_600_delayed_14_0_630_inst_req_1;
      W_send3_3_600_delayed_14_0_630_inst_ack_1<= rack(0);
      W_send3_3_600_delayed_14_0_630_inst : InterlockBuffer generic map ( -- 
        name => "W_send3_3_600_delayed_14_0_630_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send3_3_606,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send3_3_600_delayed_14_0_632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send3_4_760_delayed_14_0_802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send3_4_760_delayed_14_0_802_inst_req_0;
      W_send3_4_760_delayed_14_0_802_inst_ack_0<= wack(0);
      rreq(0) <= W_send3_4_760_delayed_14_0_802_inst_req_1;
      W_send3_4_760_delayed_14_0_802_inst_ack_1<= rack(0);
      W_send3_4_760_delayed_14_0_802_inst : InterlockBuffer generic map ( -- 
        name => "W_send3_4_760_delayed_14_0_802_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send3_4_778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send3_4_760_delayed_14_0_804,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send4_1_284_delayed_14_0_293_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send4_1_284_delayed_14_0_293_inst_req_0;
      W_send4_1_284_delayed_14_0_293_inst_ack_0<= wack(0);
      rreq(0) <= W_send4_1_284_delayed_14_0_293_inst_req_1;
      W_send4_1_284_delayed_14_0_293_inst_ack_1<= rack(0);
      W_send4_1_284_delayed_14_0_293_inst : InterlockBuffer generic map ( -- 
        name => "W_send4_1_284_delayed_14_0_293_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send4_1_271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send4_1_284_delayed_14_0_295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send4_2_444_delayed_14_0_465_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send4_2_444_delayed_14_0_465_inst_req_0;
      W_send4_2_444_delayed_14_0_465_inst_ack_0<= wack(0);
      rreq(0) <= W_send4_2_444_delayed_14_0_465_inst_req_1;
      W_send4_2_444_delayed_14_0_465_inst_ack_1<= rack(0);
      W_send4_2_444_delayed_14_0_465_inst : InterlockBuffer generic map ( -- 
        name => "W_send4_2_444_delayed_14_0_465_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send4_2_443,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send4_2_444_delayed_14_0_467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send4_3_604_delayed_14_0_637_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send4_3_604_delayed_14_0_637_inst_req_0;
      W_send4_3_604_delayed_14_0_637_inst_ack_0<= wack(0);
      rreq(0) <= W_send4_3_604_delayed_14_0_637_inst_req_1;
      W_send4_3_604_delayed_14_0_637_inst_ack_1<= rack(0);
      W_send4_3_604_delayed_14_0_637_inst : InterlockBuffer generic map ( -- 
        name => "W_send4_3_604_delayed_14_0_637_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send4_3_615,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send4_3_604_delayed_14_0_639,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send4_4_764_delayed_14_0_809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send4_4_764_delayed_14_0_809_inst_req_0;
      W_send4_4_764_delayed_14_0_809_inst_ack_0<= wack(0);
      rreq(0) <= W_send4_4_764_delayed_14_0_809_inst_req_1;
      W_send4_4_764_delayed_14_0_809_inst_ack_1<= rack(0);
      W_send4_4_764_delayed_14_0_809_inst : InterlockBuffer generic map ( -- 
        name => "W_send4_4_764_delayed_14_0_809_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send4_4_787,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send4_4_764_delayed_14_0_811,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_139_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_139_final_reg_req_0;
      addr_of_139_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_139_final_reg_req_1;
      addr_of_139_final_reg_ack_1<= rack(0);
      addr_of_139_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_139_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_138_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_312_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_312_final_reg_req_0;
      addr_of_312_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_312_final_reg_req_1;
      addr_of_312_final_reg_ack_1<= rack(0);
      addr_of_312_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_312_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_311_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_484_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_484_final_reg_req_0;
      addr_of_484_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_484_final_reg_req_1;
      addr_of_484_final_reg_ack_1<= rack(0);
      addr_of_484_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_484_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_483_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr3_485,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_656_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_656_final_reg_req_0;
      addr_of_656_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_656_final_reg_req_1;
      addr_of_656_final_reg_ack_1<= rack(0);
      addr_of_656_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_656_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_655_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr4_657,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_210_48_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_210_48_buf_req_0;
      n_address1_210_48_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_210_48_buf_req_1;
      n_address1_210_48_buf_ack_1<= rack(0);
      n_address1_210_48_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_210_48_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_210_48_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_382_51_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_382_51_buf_req_0;
      n_address2_382_51_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_382_51_buf_req_1;
      n_address2_382_51_buf_ack_1<= rack(0);
      n_address2_382_51_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_382_51_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_382_51_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address3_554_56_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address3_554_56_buf_req_0;
      n_address3_554_56_buf_ack_0<= wack(0);
      rreq(0) <= n_address3_554_56_buf_req_1;
      n_address3_554_56_buf_ack_1<= rack(0);
      n_address3_554_56_buf : InterlockBuffer generic map ( -- 
        name => "n_address3_554_56_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address3_554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address3_554_56_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address4_726_65_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address4_726_65_buf_req_0;
      n_address4_726_65_buf_ack_0<= wack(0);
      rreq(0) <= n_address4_726_65_buf_req_1;
      n_address4_726_65_buf_ack_1<= rack(0);
      n_address4_726_65_buf : InterlockBuffer generic map ( -- 
        name => "n_address4_726_65_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address4_726,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address4_726_65_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter1_185_70_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter1_185_70_buf_req_0;
      n_mycounter1_185_70_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter1_185_70_buf_req_1;
      n_mycounter1_185_70_buf_ack_1<= rack(0);
      n_mycounter1_185_70_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter1_185_70_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter1_185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter1_185_70_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter2_357_75_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter2_357_75_buf_req_0;
      n_mycounter2_357_75_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter2_357_75_buf_req_1;
      n_mycounter2_357_75_buf_ack_1<= rack(0);
      n_mycounter2_357_75_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter2_357_75_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter2_357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter2_357_75_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter3_529_80_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter3_529_80_buf_req_0;
      n_mycounter3_529_80_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter3_529_80_buf_req_1;
      n_mycounter3_529_80_buf_ack_1<= rack(0);
      n_mycounter3_529_80_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter3_529_80_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter3_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter3_529_80_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter4_701_85_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter4_701_85_buf_req_0;
      n_mycounter4_701_85_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter4_701_85_buf_req_1;
      n_mycounter4_701_85_buf_ack_1<= rack(0);
      n_mycounter4_701_85_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter4_701_85_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter4_701,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter4_701_85_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row1_193_88_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row1_193_88_buf_req_0;
      n_row1_193_88_buf_ack_0<= wack(0);
      rreq(0) <= n_row1_193_88_buf_req_1;
      n_row1_193_88_buf_ack_1<= rack(0);
      n_row1_193_88_buf : InterlockBuffer generic map ( -- 
        name => "n_row1_193_88_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row1_193,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row1_193_88_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row2_365_95_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row2_365_95_buf_req_0;
      n_row2_365_95_buf_ack_0<= wack(0);
      rreq(0) <= n_row2_365_95_buf_req_1;
      n_row2_365_95_buf_ack_1<= rack(0);
      n_row2_365_95_buf : InterlockBuffer generic map ( -- 
        name => "n_row2_365_95_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row2_365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row2_365_95_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row3_537_100_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row3_537_100_buf_req_0;
      n_row3_537_100_buf_ack_0<= wack(0);
      rreq(0) <= n_row3_537_100_buf_req_1;
      n_row3_537_100_buf_ack_1<= rack(0);
      n_row3_537_100_buf : InterlockBuffer generic map ( -- 
        name => "n_row3_537_100_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row3_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row3_537_100_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row4_709_105_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row4_709_105_buf_req_0;
      n_row4_709_105_buf_ack_0<= wack(0);
      rreq(0) <= n_row4_709_105_buf_req_1;
      n_row4_709_105_buf_ack_1<= rack(0);
      n_row4_709_105_buf : InterlockBuffer generic map ( -- 
        name => "n_row4_709_105_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row4_709,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row4_709_105_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_start1_168_110_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_start1_168_110_buf_req_0;
      n_start1_168_110_buf_ack_0<= wack(0);
      rreq(0) <= n_start1_168_110_buf_req_1;
      n_start1_168_110_buf_ack_1<= rack(0);
      n_start1_168_110_buf : InterlockBuffer generic map ( -- 
        name => "n_start1_168_110_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_start1_168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_start1_168_110_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_start2_340_115_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_start2_340_115_buf_req_0;
      n_start2_340_115_buf_ack_0<= wack(0);
      rreq(0) <= n_start2_340_115_buf_req_1;
      n_start2_340_115_buf_ack_1<= rack(0);
      n_start2_340_115_buf : InterlockBuffer generic map ( -- 
        name => "n_start2_340_115_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_start2_340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_start2_340_115_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_start3_512_120_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_start3_512_120_buf_req_0;
      n_start3_512_120_buf_ack_0<= wack(0);
      rreq(0) <= n_start3_512_120_buf_req_1;
      n_start3_512_120_buf_ack_1<= rack(0);
      n_start3_512_120_buf : InterlockBuffer generic map ( -- 
        name => "n_start3_512_120_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_start3_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_start3_512_120_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_start4_684_125_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_start4_684_125_buf_req_0;
      n_start4_684_125_buf_ack_0<= wack(0);
      rreq(0) <= n_start4_684_125_buf_req_1;
      n_start4_684_125_buf_ack_1<= rack(0);
      n_start4_684_125_buf : InterlockBuffer generic map ( -- 
        name => "n_start4_684_125_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_start4_684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_start4_684_125_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_164_inst
    process(address1_44) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := address1_44(1 downto 0);
      last2_1_165 <= tmp_var; -- 
    end process;
    -- interlock type_cast_180_inst
    process(last2_1_165) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := last2_1_165(1 downto 0);
      type_cast_180_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_200_inst
    process(ADD_u32_u32_199_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ADD_u32_u32_199_wire(31 downto 0);
      type_cast_200_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_204_inst
    process(last2_1_165) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := last2_1_165(1 downto 0);
      type_cast_204_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_336_inst
    process(address2_49) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := address2_49(1 downto 0);
      last2_2_337 <= tmp_var; -- 
    end process;
    -- interlock type_cast_352_inst
    process(last2_2_337) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := last2_2_337(1 downto 0);
      type_cast_352_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_35_inst
    process(MUL_u16_u16_34_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_34_wire(15 downto 0);
      m_factor_36 <= tmp_var; -- 
    end process;
    -- interlock type_cast_372_inst
    process(ADD_u32_u32_371_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ADD_u32_u32_371_wire(31 downto 0);
      type_cast_372_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_376_inst
    process(last2_2_337) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := last2_2_337(1 downto 0);
      type_cast_376_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_508_inst
    process(address3_54) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := address3_54(1 downto 0);
      last2_3_509 <= tmp_var; -- 
    end process;
    -- interlock type_cast_524_inst
    process(last2_3_509) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := last2_3_509(1 downto 0);
      type_cast_524_wire <= tmp_var; -- 
    end process;
    type_cast_53_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_53_inst_req_0;
      type_cast_53_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_53_inst_req_1;
      type_cast_53_inst_ack_1<= rack(0);
      type_cast_53_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_53_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_53_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_544_inst
    process(ADD_u32_u32_543_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ADD_u32_u32_543_wire(31 downto 0);
      type_cast_544_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_548_inst
    process(last2_3_509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := last2_3_509(1 downto 0);
      type_cast_548_wire <= tmp_var; -- 
    end process;
    type_cast_58_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_58_inst_req_0;
      type_cast_58_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_58_inst_req_1;
      type_cast_58_inst_ack_1<= rack(0);
      type_cast_58_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_58_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m2_factor_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_58_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u32_u32_63_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_64_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_680_inst
    process(address4_59) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := address4_59(1 downto 0);
      last2_4_681 <= tmp_var; -- 
    end process;
    -- interlock type_cast_696_inst
    process(last2_4_681) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := last2_4_681(1 downto 0);
      type_cast_696_wire <= tmp_var; -- 
    end process;
    type_cast_69_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_69_inst_req_0;
      type_cast_69_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_69_inst_req_1;
      type_cast_69_inst_ack_1<= rack(0);
      type_cast_69_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_69_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_69_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_716_inst
    process(ADD_u32_u32_715_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ADD_u32_u32_715_wire(31 downto 0);
      type_cast_716_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_720_inst
    process(last2_4_681) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := last2_4_681(1 downto 0);
      type_cast_720_wire <= tmp_var; -- 
    end process;
    type_cast_74_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_74_inst_req_0;
      type_cast_74_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_74_inst_req_1;
      type_cast_74_inst_ack_1<= rack(0);
      type_cast_74_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_74_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_74_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_79_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_79_inst_req_0;
      type_cast_79_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_79_inst_req_1;
      type_cast_79_inst_ack_1<= rack(0);
      type_cast_79_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_79_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_79_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_84_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_84_inst_req_0;
      type_cast_84_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_84_inst_req_1;
      type_cast_84_inst_ack_1<= rack(0);
      type_cast_84_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_84_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_84_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_138_index_1_rename
    process(LSHR_u64_u64_137_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_137_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_137_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_138_index_1_resize
    process(LSHR_u64_u64_137_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_137_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_137_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_138_root_address_inst
    process(array_obj_ref_138_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_138_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_138_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_311_index_1_rename
    process(LSHR_u64_u64_310_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_310_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_310_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_311_index_1_resize
    process(LSHR_u64_u64_310_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_310_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_310_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_311_root_address_inst
    process(array_obj_ref_311_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_311_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_311_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_483_index_1_rename
    process(LSHR_u64_u64_482_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_482_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_482_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_483_index_1_resize
    process(LSHR_u64_u64_482_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_482_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_482_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_483_root_address_inst
    process(array_obj_ref_483_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_483_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_483_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_655_index_1_rename
    process(LSHR_u64_u64_654_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_654_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_654_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_655_index_1_resize
    process(LSHR_u64_u64_654_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_654_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_654_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_655_root_address_inst
    process(array_obj_ref_655_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_655_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_655_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_143_addr_0
    process(ptr_deref_143_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_143_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_143_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_143_base_resize
    process(fetch_addr1_140) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_140;
      ov := iv(13 downto 0);
      ptr_deref_143_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_143_gather_scatter
    process(ptr_deref_143_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_143_data_0;
      ov(63 downto 0) := iv;
      fv1_144 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_143_root_address_inst
    process(ptr_deref_143_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_143_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_143_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_316_addr_0
    process(ptr_deref_316_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_316_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_316_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_316_base_resize
    process(fetch_addr2_313) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_313;
      ov := iv(13 downto 0);
      ptr_deref_316_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_316_gather_scatter
    process(ptr_deref_316_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_316_data_0;
      ov(63 downto 0) := iv;
      fv2_317 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_316_root_address_inst
    process(ptr_deref_316_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_316_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_316_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_addr_0
    process(ptr_deref_488_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_488_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_488_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_base_resize
    process(fetch_addr3_485) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr3_485;
      ov := iv(13 downto 0);
      ptr_deref_488_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_gather_scatter
    process(ptr_deref_488_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_488_data_0;
      ov(63 downto 0) := iv;
      fv3_489 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_root_address_inst
    process(ptr_deref_488_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_488_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_488_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_660_addr_0
    process(ptr_deref_660_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_660_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_660_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_660_base_resize
    process(fetch_addr4_657) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr4_657;
      ov := iv(13 downto 0);
      ptr_deref_660_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_660_gather_scatter
    process(ptr_deref_660_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_660_data_0;
      ov(63 downto 0) := iv;
      fv4_661 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_660_root_address_inst
    process(ptr_deref_660_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_660_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_660_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_42_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= OR_u1_u1_823_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_42_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_42_branch_req_0,
          ack0 => do_while_stmt_42_branch_ack_0,
          ack1 => do_while_stmt_42_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_190_inst
    process(row1_86) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row1_86, konst_189_wire_constant, tmp_var);
      ADD_u16_u16_190_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_362_inst
    process(row2_91) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row2_91, konst_361_wire_constant, tmp_var);
      ADD_u16_u16_362_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_534_inst
    process(row3_96) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row3_96, konst_533_wire_constant, tmp_var);
      ADD_u16_u16_534_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_706_inst
    process(row4_101) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row4_101, konst_705_wire_constant, tmp_var);
      ADD_u16_u16_706_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_181_inst
    process(tmp_cnt1_173, type_cast_180_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp_cnt1_173, type_cast_180_wire, tmp_var);
      ADD_u32_u32_181_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_199_inst
    process(m_factor_36, mycounter1_66) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, mycounter1_66, tmp_var);
      ADD_u32_u32_199_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_353_inst
    process(tmp_cnt2_345, type_cast_352_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp_cnt2_345, type_cast_352_wire, tmp_var);
      ADD_u32_u32_353_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_371_inst
    process(m_factor_36, mycounter2_71) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, mycounter2_71, tmp_var);
      ADD_u32_u32_371_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_525_inst
    process(tmp_cnt3_517, type_cast_524_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp_cnt3_517, type_cast_524_wire, tmp_var);
      ADD_u32_u32_525_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_543_inst
    process(m_factor_36, mycounter3_76) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, mycounter3_76, tmp_var);
      ADD_u32_u32_543_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_63_inst
    process(m_factor_36, m2_factor_41) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, m2_factor_41, tmp_var);
      ADD_u32_u32_63_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_697_inst
    process(tmp_cnt4_689, type_cast_696_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp_cnt4_689, type_cast_696_wire, tmp_var);
      ADD_u32_u32_697_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_715_inst
    process(m_factor_36, mycounter4_81) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, mycounter4_81, tmp_var);
      ADD_u32_u32_715_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_209_inst
    process(address1_44, MUX_208_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_44, MUX_208_wire, tmp_var);
      n_address1_210 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_381_inst
    process(address2_49, MUX_380_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_49, MUX_380_wire, tmp_var);
      n_address2_382 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_553_inst
    process(address3_54, MUX_552_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address3_54, MUX_552_wire, tmp_var);
      n_address3_554 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_725_inst
    process(address4_59, MUX_724_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address4_59, MUX_724_wire, tmp_var);
      n_address4_726 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_229_inst
    process(send_flag1_215, OR_u1_u1_228_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag1_215, OR_u1_u1_228_wire, tmp_var);
      send1_1_230 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_237_inst
    process(start1_106, ULE_u2_u1_236_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(start1_106, ULE_u2_u1_236_wire, tmp_var);
      AND_u1_u1_237_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_243_inst
    process(NOT_u1_u1_239_wire, UGT_u32_u1_242_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_239_wire, UGT_u32_u1_242_wire, tmp_var);
      AND_u1_u1_243_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_245_inst
    process(send_flag1_215, OR_u1_u1_244_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag1_215, OR_u1_u1_244_wire, tmp_var);
      send2_1_246 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_253_inst
    process(start1_106, ULE_u2_u1_252_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(start1_106, ULE_u2_u1_252_wire, tmp_var);
      AND_u1_u1_253_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_259_inst
    process(NOT_u1_u1_255_wire, UGT_u32_u1_258_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_255_wire, UGT_u32_u1_258_wire, tmp_var);
      AND_u1_u1_259_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_261_inst
    process(send_flag1_215, OR_u1_u1_260_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag1_215, OR_u1_u1_260_wire, tmp_var);
      send3_1_262 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_270_inst
    process(send_flag1_215, OR_u1_u1_269_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag1_215, OR_u1_u1_269_wire, tmp_var);
      send4_1_271 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_401_inst
    process(send_flag2_387, OR_u1_u1_400_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag2_387, OR_u1_u1_400_wire, tmp_var);
      send1_2_402 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_409_inst
    process(start2_111, ULE_u2_u1_408_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(start2_111, ULE_u2_u1_408_wire, tmp_var);
      AND_u1_u1_409_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_415_inst
    process(NOT_u1_u1_411_wire, UGT_u32_u1_414_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_411_wire, UGT_u32_u1_414_wire, tmp_var);
      AND_u1_u1_415_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_417_inst
    process(send_flag2_387, OR_u1_u1_416_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag2_387, OR_u1_u1_416_wire, tmp_var);
      send2_2_418 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_425_inst
    process(start2_111, ULE_u2_u1_424_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(start2_111, ULE_u2_u1_424_wire, tmp_var);
      AND_u1_u1_425_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_431_inst
    process(NOT_u1_u1_427_wire, UGT_u32_u1_430_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_427_wire, UGT_u32_u1_430_wire, tmp_var);
      AND_u1_u1_431_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_433_inst
    process(send_flag2_387, OR_u1_u1_432_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag2_387, OR_u1_u1_432_wire, tmp_var);
      send3_2_434 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_442_inst
    process(send_flag2_387, OR_u1_u1_441_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag2_387, OR_u1_u1_441_wire, tmp_var);
      send4_2_443 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_573_inst
    process(send_flag3_559, OR_u1_u1_572_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag3_559, OR_u1_u1_572_wire, tmp_var);
      send1_3_574 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_581_inst
    process(start3_116, ULE_u2_u1_580_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(start3_116, ULE_u2_u1_580_wire, tmp_var);
      AND_u1_u1_581_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_587_inst
    process(NOT_u1_u1_583_wire, UGT_u32_u1_586_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_583_wire, UGT_u32_u1_586_wire, tmp_var);
      AND_u1_u1_587_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_589_inst
    process(send_flag3_559, OR_u1_u1_588_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag3_559, OR_u1_u1_588_wire, tmp_var);
      send2_3_590 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_597_inst
    process(start3_116, ULE_u2_u1_596_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(start3_116, ULE_u2_u1_596_wire, tmp_var);
      AND_u1_u1_597_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_603_inst
    process(NOT_u1_u1_599_wire, UGT_u32_u1_602_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_599_wire, UGT_u32_u1_602_wire, tmp_var);
      AND_u1_u1_603_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_605_inst
    process(send_flag3_559, OR_u1_u1_604_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag3_559, OR_u1_u1_604_wire, tmp_var);
      send3_3_606 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_614_inst
    process(send_flag3_559, OR_u1_u1_613_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag3_559, OR_u1_u1_613_wire, tmp_var);
      send4_3_615 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_745_inst
    process(send_flag4_731, OR_u1_u1_744_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag4_731, OR_u1_u1_744_wire, tmp_var);
      send1_4_746 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_753_inst
    process(start4_121, ULE_u2_u1_752_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(start4_121, ULE_u2_u1_752_wire, tmp_var);
      AND_u1_u1_753_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_759_inst
    process(NOT_u1_u1_755_wire, UGT_u32_u1_758_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_755_wire, UGT_u32_u1_758_wire, tmp_var);
      AND_u1_u1_759_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_761_inst
    process(send_flag4_731, OR_u1_u1_760_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag4_731, OR_u1_u1_760_wire, tmp_var);
      send2_4_762 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_769_inst
    process(start4_121, ULE_u2_u1_768_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(start4_121, ULE_u2_u1_768_wire, tmp_var);
      AND_u1_u1_769_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_775_inst
    process(NOT_u1_u1_771_wire, UGT_u32_u1_774_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_771_wire, UGT_u32_u1_774_wire, tmp_var);
      AND_u1_u1_775_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_777_inst
    process(send_flag4_731, OR_u1_u1_776_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag4_731, OR_u1_u1_776_wire, tmp_var);
      send3_4_778 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_786_inst
    process(send_flag4_731, OR_u1_u1_785_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(send_flag4_731, OR_u1_u1_785_wire, tmp_var);
      send4_4_787 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_225_inst
    process(last2_1_165) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last2_1_165, konst_224_wire_constant, tmp_var);
      EQ_u2_u1_225_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_397_inst
    process(last2_2_337) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last2_2_337, konst_396_wire_constant, tmp_var);
      EQ_u2_u1_397_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_569_inst
    process(last2_3_509) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last2_3_509, konst_568_wire_constant, tmp_var);
      EQ_u2_u1_569_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_741_inst
    process(last2_4_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last2_4_681, konst_740_wire_constant, tmp_var);
      EQ_u2_u1_741_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_137_inst
    process(address1_44) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_44, konst_136_wire_constant, tmp_var);
      LSHR_u64_u64_137_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_310_inst
    process(address2_49) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_49, konst_309_wire_constant, tmp_var);
      LSHR_u64_u64_310_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_482_inst
    process(address3_54) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address3_54, konst_481_wire_constant, tmp_var);
      LSHR_u64_u64_482_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_654_inst
    process(address4_59) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address4_59, konst_653_wire_constant, tmp_var);
      LSHR_u64_u64_654_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_34_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_34_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_227_inst
    process(start1_106) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start1_106, tmp_var);
      NOT_u1_u1_227_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_239_inst
    process(start1_106) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start1_106, tmp_var);
      NOT_u1_u1_239_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_255_inst
    process(start1_106) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start1_106, tmp_var);
      NOT_u1_u1_255_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_399_inst
    process(start2_111) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start2_111, tmp_var);
      NOT_u1_u1_399_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_411_inst
    process(start2_111) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start2_111, tmp_var);
      NOT_u1_u1_411_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_427_inst
    process(start2_111) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start2_111, tmp_var);
      NOT_u1_u1_427_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_571_inst
    process(start3_116) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start3_116, tmp_var);
      NOT_u1_u1_571_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_583_inst
    process(start3_116) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start3_116, tmp_var);
      NOT_u1_u1_583_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_599_inst
    process(start3_116) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start3_116, tmp_var);
      NOT_u1_u1_599_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_743_inst
    process(start4_121) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start4_121, tmp_var);
      NOT_u1_u1_743_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_755_inst
    process(start4_121) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start4_121, tmp_var);
      NOT_u1_u1_755_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_771_inst
    process(start4_121) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", start4_121, tmp_var);
      NOT_u1_u1_771_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_228_inst
    process(EQ_u2_u1_225_wire, NOT_u1_u1_227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_225_wire, NOT_u1_u1_227_wire, tmp_var);
      OR_u1_u1_228_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_244_inst
    process(AND_u1_u1_237_wire, AND_u1_u1_243_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_237_wire, AND_u1_u1_243_wire, tmp_var);
      OR_u1_u1_244_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_260_inst
    process(AND_u1_u1_253_wire, AND_u1_u1_259_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_253_wire, AND_u1_u1_259_wire, tmp_var);
      OR_u1_u1_260_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_269_inst
    process(start1_106, UGT_u32_u1_268_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(start1_106, UGT_u32_u1_268_wire, tmp_var);
      OR_u1_u1_269_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_400_inst
    process(EQ_u2_u1_397_wire, NOT_u1_u1_399_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_397_wire, NOT_u1_u1_399_wire, tmp_var);
      OR_u1_u1_400_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_416_inst
    process(AND_u1_u1_409_wire, AND_u1_u1_415_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_409_wire, AND_u1_u1_415_wire, tmp_var);
      OR_u1_u1_416_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_432_inst
    process(AND_u1_u1_425_wire, AND_u1_u1_431_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_425_wire, AND_u1_u1_431_wire, tmp_var);
      OR_u1_u1_432_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_441_inst
    process(start2_111, UGT_u32_u1_440_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(start2_111, UGT_u32_u1_440_wire, tmp_var);
      OR_u1_u1_441_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_572_inst
    process(EQ_u2_u1_569_wire, NOT_u1_u1_571_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_569_wire, NOT_u1_u1_571_wire, tmp_var);
      OR_u1_u1_572_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_588_inst
    process(AND_u1_u1_581_wire, AND_u1_u1_587_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_581_wire, AND_u1_u1_587_wire, tmp_var);
      OR_u1_u1_588_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_604_inst
    process(AND_u1_u1_597_wire, AND_u1_u1_603_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_597_wire, AND_u1_u1_603_wire, tmp_var);
      OR_u1_u1_604_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_613_inst
    process(start3_116, UGT_u32_u1_612_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(start3_116, UGT_u32_u1_612_wire, tmp_var);
      OR_u1_u1_613_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_744_inst
    process(EQ_u2_u1_741_wire, NOT_u1_u1_743_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_741_wire, NOT_u1_u1_743_wire, tmp_var);
      OR_u1_u1_744_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_760_inst
    process(AND_u1_u1_753_wire, AND_u1_u1_759_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_753_wire, AND_u1_u1_759_wire, tmp_var);
      OR_u1_u1_760_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_776_inst
    process(AND_u1_u1_769_wire, AND_u1_u1_775_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_769_wire, AND_u1_u1_775_wire, tmp_var);
      OR_u1_u1_776_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_785_inst
    process(start4_121, UGT_u32_u1_784_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(start4_121, UGT_u32_u1_784_wire, tmp_var);
      OR_u1_u1_785_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_819_inst
    process(continue_flag1_220, continue_flag2_392) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(continue_flag1_220, continue_flag2_392, tmp_var);
      OR_u1_u1_819_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_822_inst
    process(continue_flag3_564, continue_flag4_736) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(continue_flag3_564, continue_flag4_736, tmp_var);
      OR_u1_u1_822_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_823_inst
    process(OR_u1_u1_819_wire, OR_u1_u1_822_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_819_wire, OR_u1_u1_822_wire, tmp_var);
      OR_u1_u1_823_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_40_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(m_factor_36, konst_39_wire_constant, tmp_var);
      m2_factor_41 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_172_inst
    process(mycounter1_66) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(mycounter1_66, konst_171_wire_constant, tmp_var);
      tmp_cnt1_173 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_344_inst
    process(mycounter2_71) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(mycounter2_71, konst_343_wire_constant, tmp_var);
      tmp_cnt2_345 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_516_inst
    process(mycounter3_76) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(mycounter3_76, konst_515_wire_constant, tmp_var);
      tmp_cnt3_517 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_688_inst
    process(mycounter4_81) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(mycounter4_81, konst_687_wire_constant, tmp_var);
      tmp_cnt4_689 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_205_inst
    process(konst_202_wire_constant, type_cast_204_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_202_wire_constant, type_cast_204_wire, tmp_var);
      SUB_u64_u64_205_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_377_inst
    process(konst_374_wire_constant, type_cast_376_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_374_wire_constant, type_cast_376_wire, tmp_var);
      SUB_u64_u64_377_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_549_inst
    process(konst_546_wire_constant, type_cast_548_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_546_wire_constant, type_cast_548_wire, tmp_var);
      SUB_u64_u64_549_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_721_inst
    process(konst_718_wire_constant, type_cast_720_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_718_wire_constant, type_cast_720_wire, tmp_var);
      SUB_u64_u64_721_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_242_inst
    process(mycounter1_66) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter1_66, konst_241_wire_constant, tmp_var);
      UGT_u32_u1_242_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_258_inst
    process(mycounter1_66) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter1_66, konst_257_wire_constant, tmp_var);
      UGT_u32_u1_258_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_268_inst
    process(mycounter1_66) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter1_66, konst_267_wire_constant, tmp_var);
      UGT_u32_u1_268_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_414_inst
    process(mycounter2_71) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter2_71, konst_413_wire_constant, tmp_var);
      UGT_u32_u1_414_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_430_inst
    process(mycounter2_71) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter2_71, konst_429_wire_constant, tmp_var);
      UGT_u32_u1_430_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_440_inst
    process(mycounter2_71) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter2_71, konst_439_wire_constant, tmp_var);
      UGT_u32_u1_440_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_586_inst
    process(mycounter3_76) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter3_76, konst_585_wire_constant, tmp_var);
      UGT_u32_u1_586_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_602_inst
    process(mycounter3_76) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter3_76, konst_601_wire_constant, tmp_var);
      UGT_u32_u1_602_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_612_inst
    process(mycounter3_76) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter3_76, konst_611_wire_constant, tmp_var);
      UGT_u32_u1_612_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_758_inst
    process(mycounter4_81) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter4_81, konst_757_wire_constant, tmp_var);
      UGT_u32_u1_758_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_774_inst
    process(mycounter4_81) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter4_81, konst_773_wire_constant, tmp_var);
      UGT_u32_u1_774_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_784_inst
    process(mycounter4_81) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mycounter4_81, konst_783_wire_constant, tmp_var);
      UGT_u32_u1_784_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u2_u1_236_inst
    process(last2_1_165) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(last2_1_165, konst_235_wire_constant, tmp_var);
      ULE_u2_u1_236_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u2_u1_252_inst
    process(last2_1_165) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(last2_1_165, konst_251_wire_constant, tmp_var);
      ULE_u2_u1_252_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u2_u1_408_inst
    process(last2_2_337) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(last2_2_337, konst_407_wire_constant, tmp_var);
      ULE_u2_u1_408_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u2_u1_424_inst
    process(last2_2_337) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(last2_2_337, konst_423_wire_constant, tmp_var);
      ULE_u2_u1_424_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u2_u1_580_inst
    process(last2_3_509) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(last2_3_509, konst_579_wire_constant, tmp_var);
      ULE_u2_u1_580_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u2_u1_596_inst
    process(last2_3_509) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(last2_3_509, konst_595_wire_constant, tmp_var);
      ULE_u2_u1_596_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u2_u1_752_inst
    process(last2_4_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(last2_4_681, konst_751_wire_constant, tmp_var);
      ULE_u2_u1_752_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u2_u1_768_inst
    process(last2_4_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(last2_4_681, konst_767_wire_constant, tmp_var);
      ULE_u2_u1_768_wire <= tmp_var; --
    end process;
    -- binary operator ULE_u32_u1_130_inst
    process(mycounter1_66) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(mycounter1_66, konst_129_wire_constant, tmp_var);
      next_row1_131 <= tmp_var; --
    end process;
    -- binary operator ULE_u32_u1_303_inst
    process(mycounter2_71) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(mycounter2_71, konst_302_wire_constant, tmp_var);
      next_row2_304 <= tmp_var; --
    end process;
    -- binary operator ULE_u32_u1_475_inst
    process(mycounter3_76) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(mycounter3_76, konst_474_wire_constant, tmp_var);
      next_row3_476 <= tmp_var; --
    end process;
    -- binary operator ULE_u32_u1_647_inst
    process(mycounter4_81) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(mycounter4_81, konst_646_wire_constant, tmp_var);
      next_row4_648 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_214_inst
    process(row1_86, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row1_86, row_in_buffer, tmp_var);
      send_flag1_215 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_219_inst
    process(n_row1_193, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row1_193, row_in_buffer, tmp_var);
      continue_flag1_220 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_386_inst
    process(row2_91, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row2_91, row_in_buffer, tmp_var);
      send_flag2_387 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_391_inst
    process(n_row2_365, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row2_365, row_in_buffer, tmp_var);
      continue_flag2_392 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_558_inst
    process(row3_96, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row3_96, row_in_buffer, tmp_var);
      send_flag3_559 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_563_inst
    process(n_row3_537, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row3_537, row_in_buffer, tmp_var);
      continue_flag3_564 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_730_inst
    process(row4_101, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row4_101, row_in_buffer, tmp_var);
      send_flag4_731 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_735_inst
    process(n_row4_709, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row4_709, row_in_buffer, tmp_var);
      continue_flag4_736 <= tmp_var; --
    end process;
    -- shared split operator group (130) : array_obj_ref_138_index_offset 
    ApIntAdd_group_130: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_137_scaled;
      array_obj_ref_138_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_138_index_offset_req_0;
      array_obj_ref_138_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_138_index_offset_req_1;
      array_obj_ref_138_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_130_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_130_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_130",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 130
    -- shared split operator group (131) : array_obj_ref_311_index_offset 
    ApIntAdd_group_131: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_310_scaled;
      array_obj_ref_311_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_311_index_offset_req_0;
      array_obj_ref_311_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_311_index_offset_req_1;
      array_obj_ref_311_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_131_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_131_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_131",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 131
    -- shared split operator group (132) : array_obj_ref_483_index_offset 
    ApIntAdd_group_132: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_482_scaled;
      array_obj_ref_483_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_483_index_offset_req_0;
      array_obj_ref_483_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_483_index_offset_req_1;
      array_obj_ref_483_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_132_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_132_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_132",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 132
    -- shared split operator group (133) : array_obj_ref_655_index_offset 
    ApIntAdd_group_133: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_654_scaled;
      array_obj_ref_655_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_655_index_offset_req_0;
      array_obj_ref_655_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_655_index_offset_req_1;
      array_obj_ref_655_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_133_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_133_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_133",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 133
    -- shared load operator group (0) : ptr_deref_143_load_0 ptr_deref_660_load_0 ptr_deref_316_load_0 ptr_deref_488_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_143_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_660_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_316_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_488_load_0_req_0;
      ptr_deref_143_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_660_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_316_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_488_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_143_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_660_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_316_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_488_load_0_req_1;
      ptr_deref_143_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_660_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_316_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_488_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 2) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 2) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_143_word_address_0 & ptr_deref_660_word_address_0 & ptr_deref_316_word_address_0 & ptr_deref_488_word_address_0;
      ptr_deref_143_data_0 <= data_out(255 downto 192);
      ptr_deref_660_data_0 <= data_out(191 downto 128);
      ptr_deref_316_data_0 <= data_out(127 downto 64);
      ptr_deref_488_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_276_inst WPIPE_input_pipe1_283_inst WPIPE_input_pipe1_290_inst WPIPE_input_pipe1_297_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_276_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_283_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_290_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_297_inst_req_0;
      WPIPE_input_pipe1_276_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_283_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_290_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_297_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_276_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_283_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_290_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_297_inst_req_1;
      WPIPE_input_pipe1_276_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_283_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_290_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_297_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send4_1_284_delayed_14_0_295(0);
      guard_vector(1)  <= send3_1_280_delayed_14_0_288(0);
      guard_vector(2)  <= send2_1_276_delayed_14_0_281(0);
      guard_vector(3)  <= send1_1_272_delayed_14_0_274(0);
      data_in <= w_11_148 & w_21_152 & w_31_156 & w_41_160;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_input_pipe2_448_inst WPIPE_input_pipe2_455_inst WPIPE_input_pipe2_462_inst WPIPE_input_pipe2_469_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe2_448_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe2_455_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe2_462_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe2_469_inst_req_0;
      WPIPE_input_pipe2_448_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe2_455_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe2_462_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe2_469_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe2_448_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe2_455_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe2_462_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe2_469_inst_req_1;
      WPIPE_input_pipe2_448_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe2_455_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe2_462_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe2_469_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send4_2_444_delayed_14_0_467(0);
      guard_vector(1)  <= send3_2_440_delayed_14_0_460(0);
      guard_vector(2)  <= send2_2_436_delayed_14_0_453(0);
      guard_vector(3)  <= send1_2_432_delayed_14_0_446(0);
      data_in <= w_12_321 & w_22_325 & w_32_329 & w_42_333;
      input_pipe2_write_1_gI: SplitGuardInterface generic map(name => "input_pipe2_write_1_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "input_pipe2", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe2_pipe_write_req(0),
          oack => input_pipe2_pipe_write_ack(0),
          odata => input_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_input_pipe3_634_inst WPIPE_input_pipe3_627_inst WPIPE_input_pipe3_620_inst WPIPE_input_pipe3_641_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe3_634_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe3_627_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe3_620_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe3_641_inst_req_0;
      WPIPE_input_pipe3_634_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe3_627_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe3_620_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe3_641_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe3_634_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe3_627_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe3_620_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe3_641_inst_req_1;
      WPIPE_input_pipe3_634_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe3_627_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe3_620_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe3_641_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send4_3_604_delayed_14_0_639(0);
      guard_vector(1)  <= send1_3_592_delayed_14_0_618(0);
      guard_vector(2)  <= send2_3_596_delayed_14_0_625(0);
      guard_vector(3)  <= send3_3_600_delayed_14_0_632(0);
      data_in <= w_33_501 & w_23_497 & w_13_493 & w_43_505;
      input_pipe3_write_2_gI: SplitGuardInterface generic map(name => "input_pipe3_write_2_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "input_pipe3", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe3_pipe_write_req(0),
          oack => input_pipe3_pipe_write_ack(0),
          odata => input_pipe3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_input_pipe4_813_inst WPIPE_input_pipe4_799_inst WPIPE_input_pipe4_806_inst WPIPE_input_pipe4_792_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe4_813_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe4_799_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe4_806_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe4_792_inst_req_0;
      WPIPE_input_pipe4_813_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe4_799_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe4_806_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe4_792_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe4_813_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe4_799_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe4_806_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe4_792_inst_req_1;
      WPIPE_input_pipe4_813_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe4_799_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe4_806_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe4_792_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send1_4_752_delayed_14_0_790(0);
      guard_vector(1)  <= send3_4_760_delayed_14_0_804(0);
      guard_vector(2)  <= send2_4_756_delayed_14_0_797(0);
      guard_vector(3)  <= send4_4_764_delayed_14_0_811(0);
      data_in <= w_44_677 & w_24_669 & w_34_673 & w_14_665;
      input_pipe4_write_3_gI: SplitGuardInterface generic map(name => "input_pipe4_write_3_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe4_write_3: OutputPortRevised -- 
        generic map ( name => "input_pipe4", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe4_pipe_write_req(0),
          oack => input_pipe4_pipe_write_ack(0),
          odata => input_pipe4_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(47 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(63 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_3789_start: Boolean;
  signal convolution3D_CP_3789_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_1885_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1509_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1509_inst_req_0 : boolean;
  signal type_cast_1513_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1496_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1496_inst_ack_0 : boolean;
  signal type_cast_1513_inst_ack_0 : boolean;
  signal type_cast_1513_inst_req_1 : boolean;
  signal type_cast_1513_inst_ack_1 : boolean;
  signal type_cast_1525_inst_req_0 : boolean;
  signal type_cast_1500_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1509_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1521_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1509_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1521_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1496_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1496_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1521_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1534_inst_req_0 : boolean;
  signal type_cast_1538_inst_ack_1 : boolean;
  signal type_cast_1538_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1546_inst_req_0 : boolean;
  signal type_cast_1538_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1534_inst_ack_0 : boolean;
  signal type_cast_1538_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1885_inst_req_1 : boolean;
  signal type_cast_1500_inst_ack_0 : boolean;
  signal type_cast_1550_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1546_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1546_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1546_inst_ack_1 : boolean;
  signal type_cast_1871_inst_ack_1 : boolean;
  signal type_cast_1525_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1903_inst_ack_0 : boolean;
  signal type_cast_1525_inst_ack_0 : boolean;
  signal type_cast_1525_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1534_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1521_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1534_inst_ack_1 : boolean;
  signal type_cast_1550_inst_req_0 : boolean;
  signal type_cast_1550_inst_ack_1 : boolean;
  signal type_cast_1500_inst_req_0 : boolean;
  signal type_cast_1550_inst_ack_0 : boolean;
  signal type_cast_1500_inst_req_1 : boolean;
  signal array_obj_ref_2130_index_offset_req_1 : boolean;
  signal type_cast_2782_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1921_inst_ack_1 : boolean;
  signal if_stmt_2091_branch_req_0 : boolean;
  signal type_cast_1925_inst_req_0 : boolean;
  signal addr_of_2131_final_reg_req_0 : boolean;
  signal addr_of_2131_final_reg_ack_0 : boolean;
  signal call_stmt_2606_call_ack_0 : boolean;
  signal addr_of_2131_final_reg_req_1 : boolean;
  signal type_cast_2630_inst_ack_0 : boolean;
  signal addr_of_2131_final_reg_ack_1 : boolean;
  signal call_stmt_2676_call_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1885_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_2709_inst_req_1 : boolean;
  signal type_cast_2630_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1903_inst_req_1 : boolean;
  signal call_stmt_2676_call_req_0 : boolean;
  signal ptr_deref_2134_store_0_req_1 : boolean;
  signal ptr_deref_2134_store_0_ack_1 : boolean;
  signal type_cast_2762_inst_ack_1 : boolean;
  signal type_cast_2792_inst_req_1 : boolean;
  signal type_cast_1925_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1885_inst_ack_0 : boolean;
  signal ptr_deref_2134_store_0_req_0 : boolean;
  signal ptr_deref_2134_store_0_ack_0 : boolean;
  signal call_stmt_2606_call_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1559_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1559_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1921_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1559_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1559_inst_ack_1 : boolean;
  signal type_cast_1563_inst_req_0 : boolean;
  signal type_cast_1563_inst_ack_0 : boolean;
  signal type_cast_1563_inst_req_1 : boolean;
  signal type_cast_1563_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1571_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1571_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1571_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1571_inst_ack_1 : boolean;
  signal type_cast_1575_inst_req_0 : boolean;
  signal type_cast_1575_inst_ack_0 : boolean;
  signal type_cast_1575_inst_req_1 : boolean;
  signal type_cast_1575_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1584_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1584_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1584_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1584_inst_ack_1 : boolean;
  signal type_cast_1588_inst_req_0 : boolean;
  signal type_cast_1588_inst_ack_0 : boolean;
  signal type_cast_1588_inst_req_1 : boolean;
  signal type_cast_1588_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1596_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1596_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1596_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1596_inst_ack_1 : boolean;
  signal type_cast_1600_inst_req_0 : boolean;
  signal type_cast_1600_inst_ack_0 : boolean;
  signal type_cast_1600_inst_req_1 : boolean;
  signal type_cast_1600_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1609_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1609_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1609_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1609_inst_ack_1 : boolean;
  signal type_cast_1613_inst_req_0 : boolean;
  signal type_cast_1613_inst_ack_0 : boolean;
  signal type_cast_1613_inst_req_1 : boolean;
  signal type_cast_1613_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1621_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1621_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1621_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1621_inst_ack_1 : boolean;
  signal type_cast_1625_inst_req_0 : boolean;
  signal type_cast_1625_inst_ack_0 : boolean;
  signal type_cast_1625_inst_req_1 : boolean;
  signal type_cast_1625_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1634_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1634_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1634_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1634_inst_ack_1 : boolean;
  signal type_cast_1638_inst_req_0 : boolean;
  signal type_cast_1638_inst_ack_0 : boolean;
  signal type_cast_1638_inst_req_1 : boolean;
  signal type_cast_1638_inst_ack_1 : boolean;
  signal type_cast_2084_inst_req_0 : boolean;
  signal ptr_deref_1951_store_0_ack_1 : boolean;
  signal if_stmt_1965_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1646_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1646_inst_ack_0 : boolean;
  signal type_cast_1889_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1646_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1646_inst_ack_1 : boolean;
  signal ptr_deref_1951_store_0_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1921_inst_ack_0 : boolean;
  signal type_cast_1650_inst_req_0 : boolean;
  signal type_cast_1943_inst_ack_1 : boolean;
  signal type_cast_1650_inst_ack_0 : boolean;
  signal type_cast_1650_inst_req_1 : boolean;
  signal type_cast_1943_inst_req_1 : boolean;
  signal type_cast_1650_inst_ack_1 : boolean;
  signal if_stmt_1965_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1659_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1659_inst_ack_0 : boolean;
  signal type_cast_1889_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1659_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1659_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1921_inst_req_0 : boolean;
  signal type_cast_1663_inst_req_0 : boolean;
  signal type_cast_1943_inst_ack_0 : boolean;
  signal type_cast_1663_inst_ack_0 : boolean;
  signal type_cast_2069_inst_ack_1 : boolean;
  signal type_cast_1663_inst_req_1 : boolean;
  signal type_cast_1943_inst_req_0 : boolean;
  signal type_cast_1663_inst_ack_1 : boolean;
  signal array_obj_ref_2130_index_offset_ack_0 : boolean;
  signal if_stmt_1965_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1671_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1671_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1671_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1671_inst_ack_1 : boolean;
  signal type_cast_2084_inst_ack_1 : boolean;
  signal type_cast_2084_inst_req_1 : boolean;
  signal ptr_deref_1951_store_0_ack_0 : boolean;
  signal type_cast_2069_inst_req_1 : boolean;
  signal type_cast_1675_inst_req_0 : boolean;
  signal type_cast_1675_inst_ack_0 : boolean;
  signal type_cast_1675_inst_req_1 : boolean;
  signal type_cast_1675_inst_ack_1 : boolean;
  signal array_obj_ref_2130_index_offset_req_0 : boolean;
  signal ptr_deref_1951_store_0_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1684_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1684_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1684_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1684_inst_ack_1 : boolean;
  signal type_cast_2084_inst_ack_0 : boolean;
  signal type_cast_1688_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1939_inst_ack_1 : boolean;
  signal type_cast_1688_inst_ack_0 : boolean;
  signal type_cast_2069_inst_ack_0 : boolean;
  signal type_cast_1688_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1939_inst_req_1 : boolean;
  signal type_cast_1688_inst_ack_1 : boolean;
  signal if_stmt_2091_branch_ack_0 : boolean;
  signal type_cast_2069_inst_req_0 : boolean;
  signal type_cast_1697_inst_req_0 : boolean;
  signal type_cast_1697_inst_ack_0 : boolean;
  signal type_cast_1697_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1939_inst_ack_0 : boolean;
  signal type_cast_1697_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1939_inst_req_0 : boolean;
  signal type_cast_1701_inst_req_0 : boolean;
  signal type_cast_1701_inst_ack_0 : boolean;
  signal type_cast_1871_inst_req_1 : boolean;
  signal type_cast_1701_inst_req_1 : boolean;
  signal type_cast_1701_inst_ack_1 : boolean;
  signal if_stmt_2091_branch_ack_1 : boolean;
  signal array_obj_ref_2130_index_offset_ack_1 : boolean;
  signal type_cast_1889_inst_ack_0 : boolean;
  signal type_cast_1907_inst_ack_1 : boolean;
  signal type_cast_1907_inst_req_1 : boolean;
  signal type_cast_1716_inst_req_0 : boolean;
  signal type_cast_1716_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2065_inst_ack_1 : boolean;
  signal type_cast_1716_inst_req_1 : boolean;
  signal type_cast_1716_inst_ack_1 : boolean;
  signal type_cast_1889_inst_req_0 : boolean;
  signal if_stmt_2016_branch_ack_0 : boolean;
  signal if_stmt_2016_branch_ack_1 : boolean;
  signal if_stmt_2016_branch_req_0 : boolean;
  signal type_cast_1907_inst_ack_0 : boolean;
  signal type_cast_1907_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2065_inst_req_1 : boolean;
  signal if_stmt_1724_branch_req_0 : boolean;
  signal if_stmt_1724_branch_ack_1 : boolean;
  signal if_stmt_1724_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1903_inst_req_0 : boolean;
  signal type_cast_1744_inst_req_0 : boolean;
  signal type_cast_1925_inst_ack_1 : boolean;
  signal type_cast_1744_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2065_inst_ack_0 : boolean;
  signal type_cast_1744_inst_req_1 : boolean;
  signal type_cast_1925_inst_req_1 : boolean;
  signal type_cast_1744_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2065_inst_req_0 : boolean;
  signal type_cast_1760_inst_req_0 : boolean;
  signal type_cast_1760_inst_ack_0 : boolean;
  signal type_cast_1760_inst_req_1 : boolean;
  signal type_cast_1760_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1903_inst_ack_1 : boolean;
  signal type_cast_1769_inst_req_0 : boolean;
  signal type_cast_1769_inst_ack_0 : boolean;
  signal type_cast_1769_inst_req_1 : boolean;
  signal type_cast_1769_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_2709_inst_ack_1 : boolean;
  signal type_cast_1779_inst_req_0 : boolean;
  signal type_cast_2630_inst_req_1 : boolean;
  signal type_cast_1779_inst_ack_0 : boolean;
  signal type_cast_1779_inst_req_1 : boolean;
  signal type_cast_2630_inst_ack_1 : boolean;
  signal type_cast_1779_inst_ack_1 : boolean;
  signal type_cast_2549_inst_req_0 : boolean;
  signal if_stmt_2556_branch_req_0 : boolean;
  signal if_stmt_2692_branch_ack_1 : boolean;
  signal array_obj_ref_1814_index_offset_req_0 : boolean;
  signal array_obj_ref_1814_index_offset_ack_0 : boolean;
  signal array_obj_ref_1814_index_offset_req_1 : boolean;
  signal array_obj_ref_1814_index_offset_ack_1 : boolean;
  signal addr_of_1815_final_reg_req_0 : boolean;
  signal ptr_deref_2599_store_0_req_0 : boolean;
  signal addr_of_1815_final_reg_ack_0 : boolean;
  signal addr_of_1815_final_reg_req_1 : boolean;
  signal addr_of_1815_final_reg_ack_1 : boolean;
  signal call_stmt_2676_call_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1818_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1818_inst_ack_0 : boolean;
  signal type_cast_2549_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1818_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1818_inst_ack_1 : boolean;
  signal call_stmt_2676_call_ack_1 : boolean;
  signal ptr_deref_2599_store_0_ack_0 : boolean;
  signal type_cast_1822_inst_req_0 : boolean;
  signal type_cast_1822_inst_ack_0 : boolean;
  signal type_cast_1822_inst_req_1 : boolean;
  signal type_cast_1822_inst_ack_1 : boolean;
  signal if_stmt_2692_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1831_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1831_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1831_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1831_inst_ack_1 : boolean;
  signal type_cast_1835_inst_req_0 : boolean;
  signal type_cast_1835_inst_ack_0 : boolean;
  signal type_cast_1835_inst_req_1 : boolean;
  signal type_cast_1835_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1849_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1849_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1849_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1849_inst_ack_1 : boolean;
  signal type_cast_1853_inst_req_0 : boolean;
  signal type_cast_1853_inst_ack_0 : boolean;
  signal type_cast_1853_inst_req_1 : boolean;
  signal type_cast_1853_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1867_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1867_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1867_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1867_inst_ack_1 : boolean;
  signal type_cast_1871_inst_req_0 : boolean;
  signal type_cast_1871_inst_ack_0 : boolean;
  signal type_cast_2141_inst_req_0 : boolean;
  signal type_cast_2141_inst_ack_0 : boolean;
  signal type_cast_2141_inst_req_1 : boolean;
  signal type_cast_2141_inst_ack_1 : boolean;
  signal type_cast_2145_inst_req_0 : boolean;
  signal type_cast_2145_inst_ack_0 : boolean;
  signal type_cast_2145_inst_req_1 : boolean;
  signal type_cast_2145_inst_ack_1 : boolean;
  signal type_cast_2149_inst_req_0 : boolean;
  signal type_cast_2149_inst_ack_0 : boolean;
  signal type_cast_2149_inst_req_1 : boolean;
  signal type_cast_2149_inst_ack_1 : boolean;
  signal if_stmt_2187_branch_req_0 : boolean;
  signal if_stmt_2187_branch_ack_1 : boolean;
  signal if_stmt_2187_branch_ack_0 : boolean;
  signal type_cast_2208_inst_req_0 : boolean;
  signal type_cast_2208_inst_ack_0 : boolean;
  signal type_cast_2208_inst_req_1 : boolean;
  signal type_cast_2208_inst_ack_1 : boolean;
  signal type_cast_2217_inst_req_0 : boolean;
  signal type_cast_2217_inst_ack_0 : boolean;
  signal type_cast_2217_inst_req_1 : boolean;
  signal type_cast_2217_inst_ack_1 : boolean;
  signal type_cast_2226_inst_req_0 : boolean;
  signal type_cast_2226_inst_ack_0 : boolean;
  signal type_cast_2226_inst_req_1 : boolean;
  signal type_cast_2226_inst_ack_1 : boolean;
  signal type_cast_2235_inst_req_0 : boolean;
  signal type_cast_2235_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2709_inst_ack_0 : boolean;
  signal type_cast_2235_inst_req_1 : boolean;
  signal type_cast_2235_inst_ack_1 : boolean;
  signal type_cast_2782_inst_ack_0 : boolean;
  signal call_stmt_2758_call_ack_0 : boolean;
  signal WPIPE_num_out_pipe_2665_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2665_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_2709_inst_req_0 : boolean;
  signal type_cast_2240_inst_req_0 : boolean;
  signal type_cast_2240_inst_ack_0 : boolean;
  signal type_cast_2240_inst_req_1 : boolean;
  signal type_cast_2240_inst_ack_1 : boolean;
  signal type_cast_2782_inst_req_0 : boolean;
  signal call_stmt_2758_call_req_0 : boolean;
  signal type_cast_2762_inst_ack_0 : boolean;
  signal type_cast_2726_inst_ack_0 : boolean;
  signal type_cast_2762_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_2665_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_2665_inst_req_0 : boolean;
  signal type_cast_2726_inst_req_0 : boolean;
  signal array_obj_ref_2275_index_offset_req_0 : boolean;
  signal array_obj_ref_2275_index_offset_ack_0 : boolean;
  signal array_obj_ref_2275_index_offset_req_1 : boolean;
  signal WPIPE_output_pipe_2613_inst_ack_1 : boolean;
  signal array_obj_ref_2275_index_offset_ack_1 : boolean;
  signal WPIPE_output_pipe_2613_inst_req_1 : boolean;
  signal addr_of_2276_final_reg_req_0 : boolean;
  signal addr_of_2276_final_reg_ack_0 : boolean;
  signal addr_of_2276_final_reg_req_1 : boolean;
  signal WPIPE_output_pipe_2613_inst_ack_0 : boolean;
  signal addr_of_2276_final_reg_ack_1 : boolean;
  signal type_cast_2792_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2279_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2613_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2279_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2279_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2279_inst_ack_1 : boolean;
  signal type_cast_2702_inst_req_0 : boolean;
  signal type_cast_2772_inst_ack_0 : boolean;
  signal type_cast_2717_inst_ack_1 : boolean;
  signal type_cast_2717_inst_req_1 : boolean;
  signal type_cast_2283_inst_req_0 : boolean;
  signal type_cast_2283_inst_ack_0 : boolean;
  signal type_cast_2283_inst_req_1 : boolean;
  signal type_cast_2283_inst_ack_1 : boolean;
  signal type_cast_2792_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2292_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2292_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2292_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2292_inst_ack_1 : boolean;
  signal type_cast_2772_inst_req_0 : boolean;
  signal type_cast_2717_inst_ack_0 : boolean;
  signal type_cast_2296_inst_req_0 : boolean;
  signal type_cast_2296_inst_ack_0 : boolean;
  signal type_cast_2296_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2610_inst_ack_1 : boolean;
  signal type_cast_2296_inst_ack_1 : boolean;
  signal type_cast_2730_inst_ack_1 : boolean;
  signal if_stmt_2692_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2310_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2610_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2310_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2310_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2310_inst_ack_1 : boolean;
  signal type_cast_2717_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_2662_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_2705_inst_ack_1 : boolean;
  signal type_cast_2314_inst_req_0 : boolean;
  signal type_cast_2314_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2705_inst_req_1 : boolean;
  signal type_cast_2314_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2610_inst_ack_0 : boolean;
  signal type_cast_2314_inst_ack_1 : boolean;
  signal type_cast_2730_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_2662_inst_req_1 : boolean;
  signal call_stmt_2758_call_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2328_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2610_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2328_inst_ack_0 : boolean;
  signal call_stmt_2758_call_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2328_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2328_inst_ack_1 : boolean;
  signal addr_of_2596_final_reg_ack_1 : boolean;
  signal addr_of_2596_final_reg_req_1 : boolean;
  signal type_cast_2332_inst_req_0 : boolean;
  signal type_cast_2332_inst_ack_0 : boolean;
  signal type_cast_2332_inst_req_1 : boolean;
  signal type_cast_2332_inst_ack_1 : boolean;
  signal type_cast_2730_inst_ack_0 : boolean;
  signal call_stmt_2680_call_ack_1 : boolean;
  signal call_stmt_2680_call_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2346_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2346_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2346_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2346_inst_ack_1 : boolean;
  signal call_stmt_2713_call_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2662_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_2662_inst_req_0 : boolean;
  signal call_stmt_2713_call_req_1 : boolean;
  signal type_cast_2350_inst_req_0 : boolean;
  signal type_cast_2350_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2705_inst_ack_0 : boolean;
  signal type_cast_2350_inst_req_1 : boolean;
  signal type_cast_2350_inst_ack_1 : boolean;
  signal type_cast_2730_inst_req_0 : boolean;
  signal call_stmt_2680_call_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2364_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2607_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2364_inst_ack_0 : boolean;
  signal if_stmt_2556_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2364_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2607_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2364_inst_ack_1 : boolean;
  signal addr_of_2596_final_reg_ack_0 : boolean;
  signal addr_of_2596_final_reg_req_0 : boolean;
  signal call_stmt_2713_call_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2705_inst_req_0 : boolean;
  signal type_cast_2368_inst_req_0 : boolean;
  signal type_cast_2368_inst_ack_0 : boolean;
  signal type_cast_2368_inst_req_1 : boolean;
  signal type_cast_2368_inst_ack_1 : boolean;
  signal call_stmt_2680_call_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2382_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2607_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2382_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2382_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2607_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2382_inst_ack_1 : boolean;
  signal call_stmt_2713_call_req_0 : boolean;
  signal type_cast_2386_inst_req_0 : boolean;
  signal type_cast_2386_inst_ack_0 : boolean;
  signal type_cast_2386_inst_req_1 : boolean;
  signal type_cast_2386_inst_ack_1 : boolean;
  signal type_cast_2772_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2400_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2400_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2400_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2400_inst_ack_1 : boolean;
  signal type_cast_2640_inst_ack_1 : boolean;
  signal type_cast_2404_inst_req_0 : boolean;
  signal type_cast_2404_inst_ack_0 : boolean;
  signal type_cast_2404_inst_req_1 : boolean;
  signal type_cast_2404_inst_ack_1 : boolean;
  signal type_cast_2772_inst_req_1 : boolean;
  signal type_cast_2782_inst_ack_1 : boolean;
  signal type_cast_2726_inst_ack_1 : boolean;
  signal type_cast_2640_inst_req_1 : boolean;
  signal type_cast_2640_inst_ack_0 : boolean;
  signal type_cast_2640_inst_req_0 : boolean;
  signal call_stmt_2606_call_ack_1 : boolean;
  signal call_stmt_2606_call_req_1 : boolean;
  signal array_obj_ref_2595_index_offset_ack_1 : boolean;
  signal array_obj_ref_2595_index_offset_req_1 : boolean;
  signal ptr_deref_2412_store_0_req_0 : boolean;
  signal ptr_deref_2412_store_0_ack_0 : boolean;
  signal ptr_deref_2412_store_0_req_1 : boolean;
  signal ptr_deref_2412_store_0_ack_1 : boolean;
  signal type_cast_2762_inst_req_1 : boolean;
  signal type_cast_2726_inst_req_1 : boolean;
  signal type_cast_2792_inst_ack_1 : boolean;
  signal array_obj_ref_2595_index_offset_ack_0 : boolean;
  signal array_obj_ref_2595_index_offset_req_0 : boolean;
  signal type_cast_2702_inst_ack_1 : boolean;
  signal type_cast_2702_inst_req_1 : boolean;
  signal if_stmt_2426_branch_req_0 : boolean;
  signal type_cast_2549_inst_ack_1 : boolean;
  signal type_cast_2549_inst_req_1 : boolean;
  signal if_stmt_2426_branch_ack_1 : boolean;
  signal ptr_deref_2599_store_0_ack_1 : boolean;
  signal if_stmt_2426_branch_ack_0 : boolean;
  signal ptr_deref_2599_store_0_req_1 : boolean;
  signal if_stmt_2556_branch_ack_1 : boolean;
  signal type_cast_2655_inst_ack_0 : boolean;
  signal type_cast_2702_inst_ack_0 : boolean;
  signal if_stmt_2477_branch_req_0 : boolean;
  signal if_stmt_2477_branch_ack_1 : boolean;
  signal if_stmt_2477_branch_ack_0 : boolean;
  signal type_cast_2492_inst_req_0 : boolean;
  signal type_cast_2492_inst_ack_0 : boolean;
  signal type_cast_2492_inst_req_1 : boolean;
  signal type_cast_2492_inst_ack_1 : boolean;
  signal type_cast_2655_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2530_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2530_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2530_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2530_inst_ack_1 : boolean;
  signal type_cast_2534_inst_req_0 : boolean;
  signal type_cast_2534_inst_ack_0 : boolean;
  signal type_cast_2534_inst_req_1 : boolean;
  signal type_cast_2534_inst_ack_1 : boolean;
  signal type_cast_2802_inst_req_0 : boolean;
  signal type_cast_2802_inst_ack_0 : boolean;
  signal type_cast_2802_inst_req_1 : boolean;
  signal type_cast_2802_inst_ack_1 : boolean;
  signal type_cast_2812_inst_req_0 : boolean;
  signal type_cast_2812_inst_ack_0 : boolean;
  signal type_cast_2812_inst_req_1 : boolean;
  signal type_cast_2812_inst_ack_1 : boolean;
  signal type_cast_2822_inst_req_0 : boolean;
  signal type_cast_2822_inst_ack_0 : boolean;
  signal type_cast_2822_inst_req_1 : boolean;
  signal type_cast_2822_inst_ack_1 : boolean;
  signal type_cast_2832_inst_req_0 : boolean;
  signal type_cast_2832_inst_ack_0 : boolean;
  signal type_cast_2832_inst_req_1 : boolean;
  signal type_cast_2832_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2834_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2834_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2834_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2834_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2837_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2837_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2837_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2837_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2840_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2840_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2840_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2840_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2843_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2843_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2843_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2843_inst_ack_1 : boolean;
  signal phi_stmt_2649_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2846_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2846_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2846_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2846_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2849_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2849_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2849_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2849_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2852_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2852_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2852_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2852_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2855_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2855_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2855_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2855_inst_ack_1 : boolean;
  signal phi_stmt_1802_req_0 : boolean;
  signal type_cast_1808_inst_req_0 : boolean;
  signal type_cast_1808_inst_ack_0 : boolean;
  signal type_cast_1808_inst_req_1 : boolean;
  signal type_cast_1808_inst_ack_1 : boolean;
  signal phi_stmt_1802_req_1 : boolean;
  signal phi_stmt_1802_ack_0 : boolean;
  signal phi_stmt_1996_req_1 : boolean;
  signal type_cast_1999_inst_req_0 : boolean;
  signal type_cast_1999_inst_ack_0 : boolean;
  signal type_cast_1999_inst_req_1 : boolean;
  signal type_cast_1999_inst_ack_1 : boolean;
  signal phi_stmt_1996_req_0 : boolean;
  signal phi_stmt_1996_ack_0 : boolean;
  signal phi_stmt_2037_req_0 : boolean;
  signal phi_stmt_2044_req_0 : boolean;
  signal type_cast_2043_inst_req_0 : boolean;
  signal type_cast_2043_inst_ack_0 : boolean;
  signal type_cast_2043_inst_req_1 : boolean;
  signal type_cast_2043_inst_ack_1 : boolean;
  signal phi_stmt_2037_req_1 : boolean;
  signal type_cast_2050_inst_req_0 : boolean;
  signal type_cast_2050_inst_ack_0 : boolean;
  signal type_cast_2050_inst_req_1 : boolean;
  signal type_cast_2050_inst_ack_1 : boolean;
  signal phi_stmt_2044_req_1 : boolean;
  signal phi_stmt_2037_ack_0 : boolean;
  signal phi_stmt_2044_ack_0 : boolean;
  signal type_cast_2101_inst_req_0 : boolean;
  signal type_cast_2101_inst_ack_0 : boolean;
  signal type_cast_2101_inst_req_1 : boolean;
  signal type_cast_2101_inst_ack_1 : boolean;
  signal phi_stmt_2098_req_0 : boolean;
  signal phi_stmt_2098_ack_0 : boolean;
  signal phi_stmt_2263_req_0 : boolean;
  signal type_cast_2269_inst_req_0 : boolean;
  signal type_cast_2269_inst_ack_0 : boolean;
  signal type_cast_2269_inst_req_1 : boolean;
  signal type_cast_2269_inst_ack_1 : boolean;
  signal phi_stmt_2263_req_1 : boolean;
  signal phi_stmt_2263_ack_0 : boolean;
  signal phi_stmt_2649_ack_0 : boolean;
  signal type_cast_2460_inst_req_0 : boolean;
  signal type_cast_2460_inst_ack_0 : boolean;
  signal type_cast_2460_inst_req_1 : boolean;
  signal type_cast_2460_inst_ack_1 : boolean;
  signal phi_stmt_2457_req_0 : boolean;
  signal phi_stmt_2457_req_1 : boolean;
  signal phi_stmt_2457_ack_0 : boolean;
  signal phi_stmt_2649_req_1 : boolean;
  signal phi_stmt_2502_req_0 : boolean;
  signal type_cast_2655_inst_ack_1 : boolean;
  signal phi_stmt_2509_req_0 : boolean;
  signal type_cast_2508_inst_req_0 : boolean;
  signal type_cast_2508_inst_ack_0 : boolean;
  signal type_cast_2508_inst_req_1 : boolean;
  signal type_cast_2508_inst_ack_1 : boolean;
  signal phi_stmt_2502_req_1 : boolean;
  signal type_cast_2655_inst_req_1 : boolean;
  signal type_cast_2515_inst_req_0 : boolean;
  signal type_cast_2515_inst_ack_0 : boolean;
  signal type_cast_2515_inst_req_1 : boolean;
  signal type_cast_2515_inst_ack_1 : boolean;
  signal phi_stmt_2509_req_1 : boolean;
  signal phi_stmt_2502_ack_0 : boolean;
  signal phi_stmt_2509_ack_0 : boolean;
  signal type_cast_2566_inst_req_0 : boolean;
  signal type_cast_2566_inst_ack_0 : boolean;
  signal type_cast_2566_inst_req_1 : boolean;
  signal type_cast_2566_inst_ack_1 : boolean;
  signal phi_stmt_2563_req_0 : boolean;
  signal phi_stmt_2563_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_3789_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_3789_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_3789_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_3789_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_3789: Block -- control-path 
    signal convolution3D_CP_3789_elements: BooleanArray(379 downto 0);
    -- 
  begin -- 
    convolution3D_CP_3789_elements(0) <= convolution3D_CP_3789_start;
    convolution3D_CP_3789_symbol <= convolution3D_CP_3789_elements(311);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1494/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/branch_block_stmt_1494__entry__
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723__entry__
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_Update/cr
      -- 
    rr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => RPIPE_maxpool_input_pipe_1496_inst_req_0); -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1513_inst_req_1); -- 
    cr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1538_inst_req_1); -- 
    cr_4040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1550_inst_req_1); -- 
    cr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1525_inst_req_1); -- 
    cr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1500_inst_req_1); -- 
    cr_4068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1563_inst_req_1); -- 
    cr_4096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1575_inst_req_1); -- 
    cr_4124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1588_inst_req_1); -- 
    cr_4152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1600_inst_req_1); -- 
    cr_4180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1613_inst_req_1); -- 
    cr_4208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1625_inst_req_1); -- 
    cr_4236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1638_inst_req_1); -- 
    cr_4264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1650_inst_req_1); -- 
    cr_4292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1663_inst_req_1); -- 
    cr_4320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1675_inst_req_1); -- 
    cr_4348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1688_inst_req_1); -- 
    cr_4362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1697_inst_req_1); -- 
    cr_4376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1701_inst_req_1); -- 
    cr_4390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(0), ack => type_cast_1716_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_update_start_
      -- 
    ra_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1496_inst_ack_0, ack => convolution3D_CP_3789_elements(1)); -- 
    cr_3914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(1), ack => RPIPE_maxpool_input_pipe_1496_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1496_update_completed_
      -- 
    ca_3915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1496_inst_ack_1, ack => convolution3D_CP_3789_elements(2)); -- 
    rr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(2), ack => type_cast_1500_inst_req_0); -- 
    rr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(2), ack => RPIPE_maxpool_input_pipe_1509_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_Sample/$exit
      -- 
    ra_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1500_inst_ack_0, ack => convolution3D_CP_3789_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1500_Update/$exit
      -- 
    ca_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1500_inst_ack_1, ack => convolution3D_CP_3789_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_Sample/$exit
      -- 
    ra_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1509_inst_ack_0, ack => convolution3D_CP_3789_elements(5)); -- 
    cr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(5), ack => RPIPE_maxpool_input_pipe_1509_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1509_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_Sample/$entry
      -- 
    ca_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1509_inst_ack_1, ack => convolution3D_CP_3789_elements(6)); -- 
    rr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(6), ack => type_cast_1513_inst_req_0); -- 
    rr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(6), ack => RPIPE_maxpool_input_pipe_1521_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_sample_completed_
      -- 
    ra_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1513_inst_ack_0, ack => convolution3D_CP_3789_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1513_update_completed_
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1513_inst_ack_1, ack => convolution3D_CP_3789_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_Update/$entry
      -- 
    ra_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1521_inst_ack_0, ack => convolution3D_CP_3789_elements(9)); -- 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(9), ack => RPIPE_maxpool_input_pipe_1521_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1521_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_sample_start_
      -- 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1521_inst_ack_1, ack => convolution3D_CP_3789_elements(10)); -- 
    rr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(10), ack => type_cast_1525_inst_req_0); -- 
    rr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(10), ack => RPIPE_maxpool_input_pipe_1534_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_Sample/$exit
      -- 
    ra_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1525_inst_ack_0, ack => convolution3D_CP_3789_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1525_Update/ca
      -- 
    ca_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1525_inst_ack_1, ack => convolution3D_CP_3789_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_Update/cr
      -- 
    ra_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1534_inst_ack_0, ack => convolution3D_CP_3789_elements(13)); -- 
    cr_3998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(13), ack => RPIPE_maxpool_input_pipe_1534_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1534_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_Sample/$entry
      -- 
    ca_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1534_inst_ack_1, ack => convolution3D_CP_3789_elements(14)); -- 
    rr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(14), ack => type_cast_1538_inst_req_0); -- 
    rr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(14), ack => RPIPE_maxpool_input_pipe_1546_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_sample_completed_
      -- 
    ra_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_0, ack => convolution3D_CP_3789_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1538_update_completed_
      -- 
    ca_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_1, ack => convolution3D_CP_3789_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_Sample/$exit
      -- 
    ra_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1546_inst_ack_0, ack => convolution3D_CP_3789_elements(17)); -- 
    cr_4026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(17), ack => RPIPE_maxpool_input_pipe_1546_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1546_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_Sample/rr
      -- 
    ca_4027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1546_inst_ack_1, ack => convolution3D_CP_3789_elements(18)); -- 
    rr_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(18), ack => type_cast_1550_inst_req_0); -- 
    rr_4049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(18), ack => RPIPE_maxpool_input_pipe_1559_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_Sample/ra
      -- 
    ra_4036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1550_inst_ack_0, ack => convolution3D_CP_3789_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1550_Update/ca
      -- 
    ca_4041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1550_inst_ack_1, ack => convolution3D_CP_3789_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_Update/cr
      -- 
    ra_4050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1559_inst_ack_0, ack => convolution3D_CP_3789_elements(21)); -- 
    cr_4054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(21), ack => RPIPE_maxpool_input_pipe_1559_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1559_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_Sample/rr
      -- 
    ca_4055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1559_inst_ack_1, ack => convolution3D_CP_3789_elements(22)); -- 
    rr_4063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(22), ack => type_cast_1563_inst_req_0); -- 
    rr_4077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(22), ack => RPIPE_maxpool_input_pipe_1571_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_Sample/ra
      -- 
    ra_4064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1563_inst_ack_0, ack => convolution3D_CP_3789_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1563_Update/ca
      -- 
    ca_4069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1563_inst_ack_1, ack => convolution3D_CP_3789_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_Update/cr
      -- 
    ra_4078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1571_inst_ack_0, ack => convolution3D_CP_3789_elements(25)); -- 
    cr_4082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(25), ack => RPIPE_maxpool_input_pipe_1571_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1571_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_Sample/rr
      -- 
    ca_4083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1571_inst_ack_1, ack => convolution3D_CP_3789_elements(26)); -- 
    rr_4091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(26), ack => type_cast_1575_inst_req_0); -- 
    rr_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(26), ack => RPIPE_maxpool_input_pipe_1584_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_Sample/ra
      -- 
    ra_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1575_inst_ack_0, ack => convolution3D_CP_3789_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1575_Update/ca
      -- 
    ca_4097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1575_inst_ack_1, ack => convolution3D_CP_3789_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_Update/cr
      -- 
    ra_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1584_inst_ack_0, ack => convolution3D_CP_3789_elements(29)); -- 
    cr_4110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(29), ack => RPIPE_maxpool_input_pipe_1584_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1584_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_Sample/rr
      -- 
    ca_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1584_inst_ack_1, ack => convolution3D_CP_3789_elements(30)); -- 
    rr_4119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(30), ack => type_cast_1588_inst_req_0); -- 
    rr_4133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(30), ack => RPIPE_maxpool_input_pipe_1596_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_Sample/ra
      -- 
    ra_4120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1588_inst_ack_0, ack => convolution3D_CP_3789_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1588_Update/ca
      -- 
    ca_4125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1588_inst_ack_1, ack => convolution3D_CP_3789_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_update_start_
      -- CP-element group 33: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_Update/cr
      -- 
    ra_4134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1596_inst_ack_0, ack => convolution3D_CP_3789_elements(33)); -- 
    cr_4138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(33), ack => RPIPE_maxpool_input_pipe_1596_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1596_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_Sample/rr
      -- 
    ca_4139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1596_inst_ack_1, ack => convolution3D_CP_3789_elements(34)); -- 
    rr_4147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(34), ack => type_cast_1600_inst_req_0); -- 
    rr_4161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(34), ack => RPIPE_maxpool_input_pipe_1609_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_Sample/ra
      -- 
    ra_4148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1600_inst_ack_0, ack => convolution3D_CP_3789_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1600_Update/ca
      -- 
    ca_4153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1600_inst_ack_1, ack => convolution3D_CP_3789_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_Update/cr
      -- 
    ra_4162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1609_inst_ack_0, ack => convolution3D_CP_3789_elements(37)); -- 
    cr_4166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(37), ack => RPIPE_maxpool_input_pipe_1609_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1609_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_Sample/rr
      -- 
    ca_4167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1609_inst_ack_1, ack => convolution3D_CP_3789_elements(38)); -- 
    rr_4189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(38), ack => RPIPE_maxpool_input_pipe_1621_inst_req_0); -- 
    rr_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(38), ack => type_cast_1613_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_Sample/ra
      -- 
    ra_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_0, ack => convolution3D_CP_3789_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1613_Update/ca
      -- 
    ca_4181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_1, ack => convolution3D_CP_3789_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_Update/cr
      -- 
    ra_4190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1621_inst_ack_0, ack => convolution3D_CP_3789_elements(41)); -- 
    cr_4194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(41), ack => RPIPE_maxpool_input_pipe_1621_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1621_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_Sample/rr
      -- 
    ca_4195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1621_inst_ack_1, ack => convolution3D_CP_3789_elements(42)); -- 
    rr_4203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(42), ack => type_cast_1625_inst_req_0); -- 
    rr_4217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(42), ack => RPIPE_maxpool_input_pipe_1634_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_Sample/ra
      -- 
    ra_4204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_0, ack => convolution3D_CP_3789_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1625_Update/ca
      -- 
    ca_4209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_1, ack => convolution3D_CP_3789_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_update_start_
      -- CP-element group 45: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_Update/cr
      -- 
    ra_4218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1634_inst_ack_0, ack => convolution3D_CP_3789_elements(45)); -- 
    cr_4222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(45), ack => RPIPE_maxpool_input_pipe_1634_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1634_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_Sample/rr
      -- 
    ca_4223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1634_inst_ack_1, ack => convolution3D_CP_3789_elements(46)); -- 
    rr_4231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(46), ack => type_cast_1638_inst_req_0); -- 
    rr_4245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(46), ack => RPIPE_maxpool_input_pipe_1646_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_Sample/ra
      -- 
    ra_4232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1638_inst_ack_0, ack => convolution3D_CP_3789_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1638_Update/ca
      -- 
    ca_4237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1638_inst_ack_1, ack => convolution3D_CP_3789_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_Update/cr
      -- 
    ra_4246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1646_inst_ack_0, ack => convolution3D_CP_3789_elements(49)); -- 
    cr_4250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(49), ack => RPIPE_maxpool_input_pipe_1646_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1646_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_Sample/rr
      -- 
    ca_4251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1646_inst_ack_1, ack => convolution3D_CP_3789_elements(50)); -- 
    rr_4259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(50), ack => type_cast_1650_inst_req_0); -- 
    rr_4273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(50), ack => RPIPE_maxpool_input_pipe_1659_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_Sample/ra
      -- 
    ra_4260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1650_inst_ack_0, ack => convolution3D_CP_3789_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1650_Update/ca
      -- 
    ca_4265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1650_inst_ack_1, ack => convolution3D_CP_3789_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_Update/cr
      -- 
    ra_4274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1659_inst_ack_0, ack => convolution3D_CP_3789_elements(53)); -- 
    cr_4278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(53), ack => RPIPE_maxpool_input_pipe_1659_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1659_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_Sample/rr
      -- 
    ca_4279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1659_inst_ack_1, ack => convolution3D_CP_3789_elements(54)); -- 
    rr_4287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(54), ack => type_cast_1663_inst_req_0); -- 
    rr_4301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(54), ack => RPIPE_maxpool_input_pipe_1671_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_Sample/ra
      -- 
    ra_4288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_0, ack => convolution3D_CP_3789_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1663_Update/ca
      -- 
    ca_4293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_1, ack => convolution3D_CP_3789_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_Update/cr
      -- 
    ra_4302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1671_inst_ack_0, ack => convolution3D_CP_3789_elements(57)); -- 
    cr_4306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(57), ack => RPIPE_maxpool_input_pipe_1671_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1671_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_Sample/rr
      -- 
    ca_4307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1671_inst_ack_1, ack => convolution3D_CP_3789_elements(58)); -- 
    rr_4315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(58), ack => type_cast_1675_inst_req_0); -- 
    rr_4329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(58), ack => RPIPE_maxpool_input_pipe_1684_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_Sample/ra
      -- 
    ra_4316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_0, ack => convolution3D_CP_3789_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1675_Update/ca
      -- 
    ca_4321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_1, ack => convolution3D_CP_3789_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_update_start_
      -- CP-element group 61: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_Update/cr
      -- 
    ra_4330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1684_inst_ack_0, ack => convolution3D_CP_3789_elements(61)); -- 
    cr_4334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(61), ack => RPIPE_maxpool_input_pipe_1684_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/RPIPE_maxpool_input_pipe_1684_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_Sample/rr
      -- 
    ca_4335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1684_inst_ack_1, ack => convolution3D_CP_3789_elements(62)); -- 
    rr_4343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(62), ack => type_cast_1688_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_Sample/ra
      -- 
    ra_4344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1688_inst_ack_0, ack => convolution3D_CP_3789_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1688_Update/ca
      -- 
    ca_4349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1688_inst_ack_1, ack => convolution3D_CP_3789_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	16 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_Sample/rr
      -- 
    rr_4357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(65), ack => type_cast_1697_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(12) & convolution3D_CP_3789_elements(16);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_Sample/ra
      -- 
    ra_4358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1697_inst_ack_0, ack => convolution3D_CP_3789_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1697_Update/ca
      -- 
    ca_4363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1697_inst_ack_1, ack => convolution3D_CP_3789_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_Sample/rr
      -- 
    rr_4371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(68), ack => type_cast_1701_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(20) & convolution3D_CP_3789_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_Sample/ra
      -- 
    ra_4372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_0, ack => convolution3D_CP_3789_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1701_Update/ca
      -- 
    ca_4377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_1, ack => convolution3D_CP_3789_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_Sample/rr
      -- 
    rr_4385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(71), ack => type_cast_1716_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(4) & convolution3D_CP_3789_elements(8) & convolution3D_CP_3789_elements(67) & convolution3D_CP_3789_elements(70);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_Sample/ra
      -- 
    ra_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1716_inst_ack_0, ack => convolution3D_CP_3789_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/type_cast_1716_Update/ca
      -- 
    ca_4391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1716_inst_ack_1, ack => convolution3D_CP_3789_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	28 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	36 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723__exit__
      -- CP-element group 74: 	 branch_block_stmt_1494/if_stmt_1724__entry__
      -- CP-element group 74: 	 branch_block_stmt_1494/assign_stmt_1497_to_assign_stmt_1723/$exit
      -- CP-element group 74: 	 branch_block_stmt_1494/if_stmt_1724_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1494/if_stmt_1724_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1494/if_stmt_1724_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1494/if_stmt_1724_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1494/R_cmp383_1725_place
      -- CP-element group 74: 	 branch_block_stmt_1494/if_stmt_1724_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1494/if_stmt_1724_else_link/$entry
      -- 
    branch_req_4399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(74), ack => if_stmt_1724_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(40) & convolution3D_CP_3789_elements(44) & convolution3D_CP_3789_elements(48) & convolution3D_CP_3789_elements(52) & convolution3D_CP_3789_elements(56) & convolution3D_CP_3789_elements(60) & convolution3D_CP_3789_elements(64) & convolution3D_CP_3789_elements(73) & convolution3D_CP_3789_elements(28) & convolution3D_CP_3789_elements(32) & convolution3D_CP_3789_elements(36);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_1494/merge_stmt_1730__exit__
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799__entry__
      -- CP-element group 75: 	 branch_block_stmt_1494/if_stmt_1724_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1494/if_stmt_1724_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1494/entry_bbx_xnph385
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1494/entry_bbx_xnph385_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/entry_bbx_xnph385_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1494/merge_stmt_1730_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1494/merge_stmt_1730_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1494/merge_stmt_1730_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1494/merge_stmt_1730_PhiAck/dummy
      -- 
    if_choice_transition_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1724_branch_ack_1, ack => convolution3D_CP_3789_elements(75)); -- 
    rr_4421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(75), ack => type_cast_1744_inst_req_0); -- 
    cr_4426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(75), ack => type_cast_1744_inst_req_1); -- 
    rr_4435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(75), ack => type_cast_1760_inst_req_0); -- 
    cr_4440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(75), ack => type_cast_1760_inst_req_1); -- 
    rr_4449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(75), ack => type_cast_1769_inst_req_0); -- 
    cr_4454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(75), ack => type_cast_1769_inst_req_1); -- 
    cr_4468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(75), ack => type_cast_1779_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	318 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_1494/if_stmt_1724_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1494/if_stmt_1724_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1494/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_1494/entry_forx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1494/entry_forx_xend_PhiReq/phi_stmt_1996/$entry
      -- CP-element group 76: 	 branch_block_stmt_1494/entry_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/$entry
      -- 
    else_choice_transition_4408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1724_branch_ack_0, ack => convolution3D_CP_3789_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_Sample/ra
      -- 
    ra_4422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1744_inst_ack_0, ack => convolution3D_CP_3789_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1744_Update/ca
      -- 
    ca_4427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1744_inst_ack_1, ack => convolution3D_CP_3789_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_Sample/ra
      -- 
    ra_4436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1760_inst_ack_0, ack => convolution3D_CP_3789_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1760_Update/ca
      -- 
    ca_4441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1760_inst_ack_1, ack => convolution3D_CP_3789_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_Sample/ra
      -- 
    ra_4450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1769_inst_ack_0, ack => convolution3D_CP_3789_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1769_Update/ca
      -- 
    ca_4455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1769_inst_ack_1, ack => convolution3D_CP_3789_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_Sample/rr
      -- 
    rr_4463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(83), ack => type_cast_1779_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(80) & convolution3D_CP_3789_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_Sample/ra
      -- 
    ra_4464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1779_inst_ack_0, ack => convolution3D_CP_3789_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/type_cast_1779_Update/ca
      -- 
    ca_4469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1779_inst_ack_1, ack => convolution3D_CP_3789_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	312 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799__exit__
      -- CP-element group 86: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_1494/assign_stmt_1735_to_assign_stmt_1799/$exit
      -- CP-element group 86: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1802/$entry
      -- CP-element group 86: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(78) & convolution3D_CP_3789_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	317 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_Sample/ack
      -- 
    ack_4498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1814_index_offset_ack_0, ack => convolution3D_CP_3789_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	317 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_request/req
      -- 
    ack_4503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1814_index_offset_ack_1, ack => convolution3D_CP_3789_elements(88)); -- 
    req_4512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(88), ack => addr_of_1815_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_request/ack
      -- 
    ack_4513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1815_final_reg_ack_0, ack => convolution3D_CP_3789_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	317 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_word_addrgen/root_register_ack
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_complete/ack
      -- 
    ack_4518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1815_final_reg_ack_1, ack => convolution3D_CP_3789_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	317 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_Update/cr
      -- 
    ra_4527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1818_inst_ack_0, ack => convolution3D_CP_3789_elements(91)); -- 
    cr_4531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(91), ack => RPIPE_maxpool_input_pipe_1818_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_Sample/rr
      -- 
    ca_4532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1818_inst_ack_1, ack => convolution3D_CP_3789_elements(92)); -- 
    rr_4540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(92), ack => type_cast_1822_inst_req_0); -- 
    rr_4554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(92), ack => RPIPE_maxpool_input_pipe_1831_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_Sample/ra
      -- 
    ra_4541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1822_inst_ack_0, ack => convolution3D_CP_3789_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	317 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_Update/ca
      -- 
    ca_4546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1822_inst_ack_1, ack => convolution3D_CP_3789_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_update_start_
      -- CP-element group 95: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_Update/cr
      -- 
    ra_4555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1831_inst_ack_0, ack => convolution3D_CP_3789_elements(95)); -- 
    cr_4559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(95), ack => RPIPE_maxpool_input_pipe_1831_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1831_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_Sample/rr
      -- 
    ca_4560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1831_inst_ack_1, ack => convolution3D_CP_3789_elements(96)); -- 
    rr_4568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(96), ack => type_cast_1835_inst_req_0); -- 
    rr_4582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(96), ack => RPIPE_maxpool_input_pipe_1849_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_Sample/ra
      -- 
    ra_4569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_0, ack => convolution3D_CP_3789_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	317 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_Update/ca
      -- 
    ca_4574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_1, ack => convolution3D_CP_3789_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_update_start_
      -- CP-element group 99: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_Update/cr
      -- 
    ra_4583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1849_inst_ack_0, ack => convolution3D_CP_3789_elements(99)); -- 
    cr_4587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(99), ack => RPIPE_maxpool_input_pipe_1849_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1849_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_Sample/rr
      -- 
    ca_4588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1849_inst_ack_1, ack => convolution3D_CP_3789_elements(100)); -- 
    rr_4596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(100), ack => type_cast_1853_inst_req_0); -- 
    rr_4610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(100), ack => RPIPE_maxpool_input_pipe_1867_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_Sample/ra
      -- 
    ra_4597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1853_inst_ack_0, ack => convolution3D_CP_3789_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	317 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_Update/ca
      -- 
    ca_4602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1853_inst_ack_1, ack => convolution3D_CP_3789_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_update_start_
      -- CP-element group 103: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_Update/cr
      -- 
    ra_4611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1867_inst_ack_0, ack => convolution3D_CP_3789_elements(103)); -- 
    cr_4615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(103), ack => RPIPE_maxpool_input_pipe_1867_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1867_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_Sample/rr
      -- 
    ca_4616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1867_inst_ack_1, ack => convolution3D_CP_3789_elements(104)); -- 
    rr_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(104), ack => type_cast_1871_inst_req_0); -- 
    rr_4638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(104), ack => RPIPE_maxpool_input_pipe_1885_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_Sample/ra
      -- 
    ra_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1871_inst_ack_0, ack => convolution3D_CP_3789_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	317 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_update_completed_
      -- 
    ca_4630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1871_inst_ack_1, ack => convolution3D_CP_3789_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_Update/cr
      -- CP-element group 107: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_update_start_
      -- CP-element group 107: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_Sample/ra
      -- 
    ra_4639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1885_inst_ack_0, ack => convolution3D_CP_3789_elements(107)); -- 
    cr_4643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(107), ack => RPIPE_maxpool_input_pipe_1885_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1885_Update/$exit
      -- 
    ca_4644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1885_inst_ack_1, ack => convolution3D_CP_3789_elements(108)); -- 
    rr_4652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(108), ack => type_cast_1889_inst_req_0); -- 
    rr_4666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(108), ack => RPIPE_maxpool_input_pipe_1903_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_sample_completed_
      -- 
    ra_4653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1889_inst_ack_0, ack => convolution3D_CP_3789_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	317 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_update_completed_
      -- 
    ca_4658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1889_inst_ack_1, ack => convolution3D_CP_3789_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_Sample/$exit
      -- 
    ra_4667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1903_inst_ack_0, ack => convolution3D_CP_3789_elements(111)); -- 
    cr_4671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(111), ack => RPIPE_maxpool_input_pipe_1903_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1903_Update/ca
      -- 
    ca_4672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1903_inst_ack_1, ack => convolution3D_CP_3789_elements(112)); -- 
    rr_4680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(112), ack => type_cast_1907_inst_req_0); -- 
    rr_4694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(112), ack => RPIPE_maxpool_input_pipe_1921_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_sample_completed_
      -- 
    ra_4681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_0, ack => convolution3D_CP_3789_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	317 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_update_completed_
      -- 
    ca_4686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_1, ack => convolution3D_CP_3789_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_update_start_
      -- CP-element group 115: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_sample_completed_
      -- 
    ra_4695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1921_inst_ack_0, ack => convolution3D_CP_3789_elements(115)); -- 
    cr_4699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(115), ack => RPIPE_maxpool_input_pipe_1921_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	119 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1921_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_sample_start_
      -- 
    ca_4700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1921_inst_ack_1, ack => convolution3D_CP_3789_elements(116)); -- 
    rr_4708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(116), ack => type_cast_1925_inst_req_0); -- 
    rr_4722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(116), ack => RPIPE_maxpool_input_pipe_1939_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_sample_completed_
      -- 
    ra_4709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1925_inst_ack_0, ack => convolution3D_CP_3789_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	317 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_Update/ca
      -- CP-element group 118: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_Update/$exit
      -- 
    ca_4714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1925_inst_ack_1, ack => convolution3D_CP_3789_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_update_start_
      -- CP-element group 119: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_sample_completed_
      -- 
    ra_4723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1939_inst_ack_0, ack => convolution3D_CP_3789_elements(119)); -- 
    cr_4727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(119), ack => RPIPE_maxpool_input_pipe_1939_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1939_update_completed_
      -- 
    ca_4728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1939_inst_ack_1, ack => convolution3D_CP_3789_elements(120)); -- 
    rr_4736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(120), ack => type_cast_1943_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_Sample/ra
      -- CP-element group 121: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_sample_completed_
      -- 
    ra_4737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1943_inst_ack_0, ack => convolution3D_CP_3789_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	317 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_Update/ca
      -- CP-element group 122: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_update_completed_
      -- 
    ca_4742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1943_inst_ack_1, ack => convolution3D_CP_3789_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: 	106 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	118 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/word_access_start/word_0/rr
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/ptr_deref_1951_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/ptr_deref_1951_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/ptr_deref_1951_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/ptr_deref_1951_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/$entry
      -- 
    rr_4780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(123), ack => ptr_deref_1951_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(122) & convolution3D_CP_3789_elements(90) & convolution3D_CP_3789_elements(94) & convolution3D_CP_3789_elements(98) & convolution3D_CP_3789_elements(102) & convolution3D_CP_3789_elements(106) & convolution3D_CP_3789_elements(110) & convolution3D_CP_3789_elements(114) & convolution3D_CP_3789_elements(118);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/word_access_start/word_0/ra
      -- CP-element group 124: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Sample/$exit
      -- 
    ra_4781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1951_store_0_ack_0, ack => convolution3D_CP_3789_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	317 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Update/word_access_complete/word_0/ca
      -- CP-element group 125: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Update/$exit
      -- 
    ca_4792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1951_store_0_ack_1, ack => convolution3D_CP_3789_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: 	87 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964__exit__
      -- CP-element group 126: 	 branch_block_stmt_1494/if_stmt_1965__entry__
      -- CP-element group 126: 	 branch_block_stmt_1494/if_stmt_1965_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_1494/if_stmt_1965_else_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_1494/if_stmt_1965_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_1494/if_stmt_1965_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_1494/if_stmt_1965_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_1494/if_stmt_1965_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_1494/R_exitcond28_1966_place
      -- CP-element group 126: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/$exit
      -- 
    branch_req_4800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(126), ack => if_stmt_1965_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(125) & convolution3D_CP_3789_elements(87);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	319 
    -- CP-element group 127: 	320 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_1494/merge_stmt_1971__exit__
      -- CP-element group 127: 	 branch_block_stmt_1494/assign_stmt_1978_to_assign_stmt_1993__entry__
      -- CP-element group 127: 	 branch_block_stmt_1494/assign_stmt_1978_to_assign_stmt_1993__exit__
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_1494/assign_stmt_1978_to_assign_stmt_1993/$exit
      -- CP-element group 127: 	 branch_block_stmt_1494/assign_stmt_1978_to_assign_stmt_1993/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/if_stmt_1965_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_1494/if_stmt_1965_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_1494/merge_stmt_1971_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_1494/merge_stmt_1971_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/merge_stmt_1971_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_1494/merge_stmt_1971_PhiAck/dummy
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1965_branch_ack_1, ack => convolution3D_CP_3789_elements(127)); -- 
    rr_6298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(127), ack => type_cast_1999_inst_req_0); -- 
    cr_6303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(127), ack => type_cast_1999_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	313 
    -- CP-element group 128: 	314 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_1494/if_stmt_1965_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_1494/if_stmt_1965_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/$entry
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/$entry
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1965_branch_ack_0, ack => convolution3D_CP_3789_elements(128)); -- 
    rr_6244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(128), ack => type_cast_1808_inst_req_0); -- 
    cr_6249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(128), ack => type_cast_1808_inst_req_1); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	323 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	342 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_1494/if_stmt_2016_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_1494/if_stmt_2016_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_1494/forx_xend_ifx_xend
      -- CP-element group 129: 	 branch_block_stmt_1494/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_1494/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_4830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2016_branch_ack_1, ack => convolution3D_CP_3789_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	323 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	324 
    -- CP-element group 130: 	325 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_1494/merge_stmt_2022__exit__
      -- CP-element group 130: 	 branch_block_stmt_1494/assign_stmt_2028_to_assign_stmt_2034__entry__
      -- CP-element group 130: 	 branch_block_stmt_1494/assign_stmt_2028_to_assign_stmt_2034__exit__
      -- CP-element group 130: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_1494/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_1494/assign_stmt_2028_to_assign_stmt_2034/$exit
      -- CP-element group 130: 	 branch_block_stmt_1494/assign_stmt_2028_to_assign_stmt_2034/$entry
      -- CP-element group 130: 	 branch_block_stmt_1494/if_stmt_2016_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_1494/if_stmt_2016_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_1494/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_1494/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_1494/merge_stmt_2022_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_1494/merge_stmt_2022_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_1494/merge_stmt_2022_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_1494/merge_stmt_2022_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/$entry
      -- CP-element group 130: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/$entry
      -- CP-element group 130: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/$entry
      -- 
    else_choice_transition_4834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2016_branch_ack_0, ack => convolution3D_CP_3789_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	337 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_update_start_
      -- CP-element group 131: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_Sample/$exit
      -- 
    ra_4851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2065_inst_ack_0, ack => convolution3D_CP_3789_elements(131)); -- 
    cr_4855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(131), ack => RPIPE_maxpool_input_pipe_2065_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_Update/$exit
      -- 
    ca_4856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2065_inst_ack_1, ack => convolution3D_CP_3789_elements(132)); -- 
    rr_4864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(132), ack => type_cast_2069_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_sample_completed_
      -- 
    ra_4865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2069_inst_ack_0, ack => convolution3D_CP_3789_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	337 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_update_completed_
      -- 
    ca_4870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2069_inst_ack_1, ack => convolution3D_CP_3789_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	337 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_Sample/ra
      -- 
    ra_4879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2084_inst_ack_0, ack => convolution3D_CP_3789_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	337 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_Update/$exit
      -- 
    ca_4884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2084_inst_ack_1, ack => convolution3D_CP_3789_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090__exit__
      -- CP-element group 137: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/$exit
      -- CP-element group 137: 	 branch_block_stmt_1494/if_stmt_2091__entry__
      -- CP-element group 137: 	 branch_block_stmt_1494/R_cmpx_xi_2092_place
      -- CP-element group 137: 	 branch_block_stmt_1494/if_stmt_2091_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_1494/if_stmt_2091_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_1494/if_stmt_2091_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_1494/if_stmt_2091_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_1494/if_stmt_2091_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_1494/if_stmt_2091_else_link/$entry
      -- 
    branch_req_4892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(137), ack => if_stmt_2091_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(134) & convolution3D_CP_3789_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	327 
    -- CP-element group 138: 	328 
    -- CP-element group 138: 	330 
    -- CP-element group 138: 	331 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_1494/if_stmt_2091_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_1494/if_stmt_2091_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2091_branch_ack_1, ack => convolution3D_CP_3789_elements(138)); -- 
    rr_6360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(138), ack => type_cast_2043_inst_req_0); -- 
    cr_6365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(138), ack => type_cast_2043_inst_req_1); -- 
    rr_6383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(138), ack => type_cast_2050_inst_req_0); -- 
    cr_6388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(138), ack => type_cast_2050_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	339 
    -- CP-element group 139: 	338 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_1494/if_stmt_2091_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_1494/if_stmt_2091_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/$entry
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/$entry
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2091_branch_ack_0, ack => convolution3D_CP_3789_elements(139)); -- 
    rr_6419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(139), ack => type_cast_2101_inst_req_0); -- 
    cr_6424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(139), ack => type_cast_2101_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	341 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_sample_complete
      -- CP-element group 140: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_Sample/ack
      -- CP-element group 140: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_Sample/$exit
      -- 
    ack_4932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2130_index_offset_ack_0, ack => convolution3D_CP_3789_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	341 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_request/req
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_Update/ack
      -- 
    ack_4937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2130_index_offset_ack_1, ack => convolution3D_CP_3789_elements(141)); -- 
    req_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(141), ack => addr_of_2131_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_request/ack
      -- CP-element group 142: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_request/$exit
      -- CP-element group 142: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_sample_completed_
      -- 
    ack_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2131_final_reg_ack_0, ack => convolution3D_CP_3789_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	341 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_word_addrgen/root_register_ack
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/ptr_deref_2134_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/ptr_deref_2134_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/ptr_deref_2134_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/ptr_deref_2134_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/word_access_start/word_0/rr
      -- CP-element group 143: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_update_completed_
      -- 
    ack_4952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2131_final_reg_ack_1, ack => convolution3D_CP_3789_elements(143)); -- 
    rr_4990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(143), ack => ptr_deref_2134_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Sample/word_access_start/word_0/ra
      -- 
    ra_4991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2134_store_0_ack_0, ack => convolution3D_CP_3789_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	341 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Update/word_access_complete/word_0/ca
      -- CP-element group 145: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_update_completed_
      -- 
    ca_5002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2134_store_0_ack_1, ack => convolution3D_CP_3789_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: 	140 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	342 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_1494/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136__exit__
      -- CP-element group 146: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/$exit
      -- CP-element group 146: 	 branch_block_stmt_1494/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_1494/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(145) & convolution3D_CP_3789_elements(140);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	342 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_Sample/ra
      -- 
    ra_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2141_inst_ack_0, ack => convolution3D_CP_3789_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	342 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_Update/ca
      -- 
    ca_5019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2141_inst_ack_1, ack => convolution3D_CP_3789_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	342 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_Sample/ra
      -- 
    ra_5028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2145_inst_ack_0, ack => convolution3D_CP_3789_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	342 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_Update/ca
      -- 
    ca_5033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2145_inst_ack_1, ack => convolution3D_CP_3789_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	342 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_Sample/ra
      -- 
    ra_5042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2149_inst_ack_0, ack => convolution3D_CP_3789_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	342 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_Update/ca
      -- 
    ca_5047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2149_inst_ack_1, ack => convolution3D_CP_3789_elements(152)); -- 
    -- CP-element group 153:  branch  join  transition  place  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (10) 
      -- CP-element group 153: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186__exit__
      -- CP-element group 153: 	 branch_block_stmt_1494/if_stmt_2187__entry__
      -- CP-element group 153: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/$exit
      -- CP-element group 153: 	 branch_block_stmt_1494/if_stmt_2187_dead_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_1494/if_stmt_2187_eval_test/$entry
      -- CP-element group 153: 	 branch_block_stmt_1494/if_stmt_2187_eval_test/$exit
      -- CP-element group 153: 	 branch_block_stmt_1494/if_stmt_2187_eval_test/branch_req
      -- CP-element group 153: 	 branch_block_stmt_1494/R_cmp161379_2188_place
      -- CP-element group 153: 	 branch_block_stmt_1494/if_stmt_2187_if_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_1494/if_stmt_2187_else_link/$entry
      -- 
    branch_req_5055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(153), ack => if_stmt_2187_branch_req_0); -- 
    convolution3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(148) & convolution3D_CP_3789_elements(150) & convolution3D_CP_3789_elements(152);
      gj_convolution3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: 	157 
    -- CP-element group 154: 	158 
    -- CP-element group 154: 	159 
    -- CP-element group 154: 	160 
    -- CP-element group 154: 	161 
    -- CP-element group 154: 	164 
    -- CP-element group 154: 	166 
    -- CP-element group 154:  members (36) 
      -- CP-element group 154: 	 branch_block_stmt_1494/merge_stmt_2193__exit__
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260__entry__
      -- CP-element group 154: 	 branch_block_stmt_1494/if_stmt_2187_if_link/$exit
      -- CP-element group 154: 	 branch_block_stmt_1494/if_stmt_2187_if_link/if_choice_transition
      -- CP-element group 154: 	 branch_block_stmt_1494/ifx_xend_bbx_xnph
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1494/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 154: 	 branch_block_stmt_1494/merge_stmt_2193_PhiReqMerge
      -- CP-element group 154: 	 branch_block_stmt_1494/merge_stmt_2193_PhiAck/$entry
      -- CP-element group 154: 	 branch_block_stmt_1494/merge_stmt_2193_PhiAck/$exit
      -- CP-element group 154: 	 branch_block_stmt_1494/merge_stmt_2193_PhiAck/dummy
      -- 
    if_choice_transition_5060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2187_branch_ack_1, ack => convolution3D_CP_3789_elements(154)); -- 
    rr_5077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(154), ack => type_cast_2208_inst_req_0); -- 
    cr_5082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(154), ack => type_cast_2208_inst_req_1); -- 
    rr_5091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(154), ack => type_cast_2217_inst_req_0); -- 
    cr_5096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(154), ack => type_cast_2217_inst_req_1); -- 
    rr_5105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(154), ack => type_cast_2226_inst_req_0); -- 
    cr_5110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(154), ack => type_cast_2226_inst_req_1); -- 
    cr_5124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(154), ack => type_cast_2235_inst_req_1); -- 
    cr_5138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(154), ack => type_cast_2240_inst_req_1); -- 
    -- CP-element group 155:  transition  place  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	352 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1494/if_stmt_2187_else_link/$exit
      -- CP-element group 155: 	 branch_block_stmt_1494/if_stmt_2187_else_link/else_choice_transition
      -- CP-element group 155: 	 branch_block_stmt_1494/ifx_xend_forx_xend215
      -- CP-element group 155: 	 branch_block_stmt_1494/ifx_xend_forx_xend215_PhiReq/$entry
      -- CP-element group 155: 	 branch_block_stmt_1494/ifx_xend_forx_xend215_PhiReq/phi_stmt_2457/$entry
      -- CP-element group 155: 	 branch_block_stmt_1494/ifx_xend_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/$entry
      -- 
    else_choice_transition_5064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2187_branch_ack_0, ack => convolution3D_CP_3789_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_Sample/ra
      -- 
    ra_5078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2208_inst_ack_0, ack => convolution3D_CP_3789_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2208_Update/ca
      -- 
    ca_5083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2208_inst_ack_1, ack => convolution3D_CP_3789_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	154 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_Sample/ra
      -- 
    ra_5092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2217_inst_ack_0, ack => convolution3D_CP_3789_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	154 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	162 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2217_Update/ca
      -- 
    ca_5097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2217_inst_ack_1, ack => convolution3D_CP_3789_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	154 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_Sample/ra
      -- 
    ra_5106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2226_inst_ack_0, ack => convolution3D_CP_3789_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	154 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2226_Update/ca
      -- 
    ca_5111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2226_inst_ack_1, ack => convolution3D_CP_3789_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	157 
    -- CP-element group 162: 	159 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_Sample/rr
      -- 
    rr_5119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(162), ack => type_cast_2235_inst_req_0); -- 
    convolution3D_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(157) & convolution3D_CP_3789_elements(159) & convolution3D_CP_3789_elements(161);
      gj_convolution3D_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_Sample/ra
      -- 
    ra_5120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2235_inst_ack_0, ack => convolution3D_CP_3789_elements(163)); -- 
    -- CP-element group 164:  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	154 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2235_Update/ca
      -- CP-element group 164: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_Sample/rr
      -- 
    ca_5125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2235_inst_ack_1, ack => convolution3D_CP_3789_elements(164)); -- 
    rr_5133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(164), ack => type_cast_2240_inst_req_0); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_Sample/ra
      -- 
    ra_5134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2240_inst_ack_0, ack => convolution3D_CP_3789_elements(165)); -- 
    -- CP-element group 166:  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	154 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	343 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260__exit__
      -- CP-element group 166: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163
      -- CP-element group 166: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/$exit
      -- CP-element group 166: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_1494/assign_stmt_2199_to_assign_stmt_2260/type_cast_2240_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_2263/$entry
      -- CP-element group 166: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/$entry
      -- 
    ca_5139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2240_inst_ack_1, ack => convolution3D_CP_3789_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	348 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	206 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_sample_complete
      -- CP-element group 167: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_Sample/ack
      -- 
    ack_5168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2275_index_offset_ack_0, ack => convolution3D_CP_3789_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	348 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (11) 
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_root_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_offset_calculated
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_Update/ack
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_base_plus_offset/$entry
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_base_plus_offset/$exit
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_request/$entry
      -- CP-element group 168: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_request/req
      -- 
    ack_5173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2275_index_offset_ack_1, ack => convolution3D_CP_3789_elements(168)); -- 
    req_5182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(168), ack => addr_of_2276_final_reg_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_request/$exit
      -- CP-element group 169: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_request/ack
      -- 
    ack_5183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2276_final_reg_ack_0, ack => convolution3D_CP_3789_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	348 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	203 
    -- CP-element group 170:  members (19) 
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_complete/$exit
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_complete/ack
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_word_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_address_resized
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_addr_resize/$entry
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_addr_resize/$exit
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_addr_resize/base_resize_req
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_addr_resize/base_resize_ack
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_word_addrgen/$entry
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_word_addrgen/$exit
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_word_addrgen/root_register_req
      -- CP-element group 170: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_word_addrgen/root_register_ack
      -- 
    ack_5188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2276_final_reg_ack_1, ack => convolution3D_CP_3789_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	348 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_update_start_
      -- CP-element group 171: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_Sample/ra
      -- CP-element group 171: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_Update/cr
      -- 
    ra_5197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2279_inst_ack_0, ack => convolution3D_CP_3789_elements(171)); -- 
    cr_5201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(171), ack => RPIPE_maxpool_input_pipe_2279_inst_req_1); -- 
    -- CP-element group 172:  fork  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: 	175 
    -- CP-element group 172:  members (9) 
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_Update/ca
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_Sample/rr
      -- 
    ca_5202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2279_inst_ack_1, ack => convolution3D_CP_3789_elements(172)); -- 
    rr_5210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(172), ack => type_cast_2283_inst_req_0); -- 
    rr_5224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(172), ack => RPIPE_maxpool_input_pipe_2292_inst_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_Sample/ra
      -- 
    ra_5211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2283_inst_ack_0, ack => convolution3D_CP_3789_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	348 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	203 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_Update/ca
      -- 
    ca_5216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2283_inst_ack_1, ack => convolution3D_CP_3789_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	172 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_Update/cr
      -- 
    ra_5225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2292_inst_ack_0, ack => convolution3D_CP_3789_elements(175)); -- 
    cr_5229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(175), ack => RPIPE_maxpool_input_pipe_2292_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2292_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_Sample/rr
      -- 
    ca_5230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2292_inst_ack_1, ack => convolution3D_CP_3789_elements(176)); -- 
    rr_5238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(176), ack => type_cast_2296_inst_req_0); -- 
    rr_5252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(176), ack => RPIPE_maxpool_input_pipe_2310_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_Sample/ra
      -- 
    ra_5239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2296_inst_ack_0, ack => convolution3D_CP_3789_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	348 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	203 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_Update/ca
      -- 
    ca_5244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2296_inst_ack_1, ack => convolution3D_CP_3789_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_update_start_
      -- CP-element group 179: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_Update/cr
      -- 
    ra_5253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2310_inst_ack_0, ack => convolution3D_CP_3789_elements(179)); -- 
    cr_5257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(179), ack => RPIPE_maxpool_input_pipe_2310_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2310_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_Sample/rr
      -- 
    ca_5258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2310_inst_ack_1, ack => convolution3D_CP_3789_elements(180)); -- 
    rr_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(180), ack => type_cast_2314_inst_req_0); -- 
    rr_5280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(180), ack => RPIPE_maxpool_input_pipe_2328_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_Sample/ra
      -- 
    ra_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2314_inst_ack_0, ack => convolution3D_CP_3789_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	348 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	203 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_Update/ca
      -- 
    ca_5272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2314_inst_ack_1, ack => convolution3D_CP_3789_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_update_start_
      -- CP-element group 183: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_Update/cr
      -- 
    ra_5281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2328_inst_ack_0, ack => convolution3D_CP_3789_elements(183)); -- 
    cr_5285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(183), ack => RPIPE_maxpool_input_pipe_2328_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2328_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_Sample/rr
      -- 
    ca_5286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2328_inst_ack_1, ack => convolution3D_CP_3789_elements(184)); -- 
    rr_5294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(184), ack => type_cast_2332_inst_req_0); -- 
    rr_5308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(184), ack => RPIPE_maxpool_input_pipe_2346_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_Sample/ra
      -- 
    ra_5295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2332_inst_ack_0, ack => convolution3D_CP_3789_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	348 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	203 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_Update/ca
      -- 
    ca_5300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2332_inst_ack_1, ack => convolution3D_CP_3789_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_update_start_
      -- CP-element group 187: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_Update/cr
      -- 
    ra_5309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2346_inst_ack_0, ack => convolution3D_CP_3789_elements(187)); -- 
    cr_5313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(187), ack => RPIPE_maxpool_input_pipe_2346_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2346_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_Sample/rr
      -- 
    ca_5314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2346_inst_ack_1, ack => convolution3D_CP_3789_elements(188)); -- 
    rr_5322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(188), ack => type_cast_2350_inst_req_0); -- 
    rr_5336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(188), ack => RPIPE_maxpool_input_pipe_2364_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_Sample/ra
      -- 
    ra_5323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2350_inst_ack_0, ack => convolution3D_CP_3789_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	348 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	203 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_Update/ca
      -- 
    ca_5328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2350_inst_ack_1, ack => convolution3D_CP_3789_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_update_start_
      -- CP-element group 191: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_Update/cr
      -- 
    ra_5337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2364_inst_ack_0, ack => convolution3D_CP_3789_elements(191)); -- 
    cr_5341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(191), ack => RPIPE_maxpool_input_pipe_2364_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2364_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_Sample/rr
      -- 
    ca_5342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2364_inst_ack_1, ack => convolution3D_CP_3789_elements(192)); -- 
    rr_5350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(192), ack => type_cast_2368_inst_req_0); -- 
    rr_5364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(192), ack => RPIPE_maxpool_input_pipe_2382_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_Sample/ra
      -- 
    ra_5351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2368_inst_ack_0, ack => convolution3D_CP_3789_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	348 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	203 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_Update/ca
      -- 
    ca_5356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2368_inst_ack_1, ack => convolution3D_CP_3789_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_update_start_
      -- CP-element group 195: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_Update/cr
      -- 
    ra_5365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2382_inst_ack_0, ack => convolution3D_CP_3789_elements(195)); -- 
    cr_5369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(195), ack => RPIPE_maxpool_input_pipe_2382_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	199 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2382_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_Sample/rr
      -- 
    ca_5370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2382_inst_ack_1, ack => convolution3D_CP_3789_elements(196)); -- 
    rr_5378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(196), ack => type_cast_2386_inst_req_0); -- 
    rr_5392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(196), ack => RPIPE_maxpool_input_pipe_2400_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_Sample/ra
      -- 
    ra_5379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2386_inst_ack_0, ack => convolution3D_CP_3789_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	348 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	203 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_Update/ca
      -- 
    ca_5384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2386_inst_ack_1, ack => convolution3D_CP_3789_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_update_start_
      -- CP-element group 199: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_Update/cr
      -- 
    ra_5393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2400_inst_ack_0, ack => convolution3D_CP_3789_elements(199)); -- 
    cr_5397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(199), ack => RPIPE_maxpool_input_pipe_2400_inst_req_1); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2400_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_Sample/rr
      -- 
    ca_5398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2400_inst_ack_1, ack => convolution3D_CP_3789_elements(200)); -- 
    rr_5406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(200), ack => type_cast_2404_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_Sample/ra
      -- 
    ra_5407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_0, ack => convolution3D_CP_3789_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	348 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_Update/ca
      -- 
    ca_5412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_1, ack => convolution3D_CP_3789_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: 	170 
    -- CP-element group 203: 	174 
    -- CP-element group 203: 	178 
    -- CP-element group 203: 	182 
    -- CP-element group 203: 	186 
    -- CP-element group 203: 	190 
    -- CP-element group 203: 	194 
    -- CP-element group 203: 	198 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (9) 
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/ptr_deref_2412_Split/$entry
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/ptr_deref_2412_Split/$exit
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/ptr_deref_2412_Split/split_req
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/ptr_deref_2412_Split/split_ack
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/word_access_start/$entry
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/word_access_start/word_0/$entry
      -- CP-element group 203: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/word_access_start/word_0/rr
      -- 
    rr_5450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(203), ack => ptr_deref_2412_store_0_req_0); -- 
    convolution3D_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(202) & convolution3D_CP_3789_elements(170) & convolution3D_CP_3789_elements(174) & convolution3D_CP_3789_elements(178) & convolution3D_CP_3789_elements(182) & convolution3D_CP_3789_elements(186) & convolution3D_CP_3789_elements(190) & convolution3D_CP_3789_elements(194) & convolution3D_CP_3789_elements(198);
      gj_convolution3D_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/word_access_start/$exit
      -- CP-element group 204: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/word_access_start/word_0/$exit
      -- CP-element group 204: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Sample/word_access_start/word_0/ra
      -- 
    ra_5451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2412_store_0_ack_0, ack => convolution3D_CP_3789_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	348 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Update/word_access_complete/$exit
      -- CP-element group 205: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Update/word_access_complete/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Update/word_access_complete/word_0/ca
      -- 
    ca_5462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2412_store_0_ack_1, ack => convolution3D_CP_3789_elements(205)); -- 
    -- CP-element group 206:  branch  join  transition  place  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	167 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (10) 
      -- CP-element group 206: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425__exit__
      -- CP-element group 206: 	 branch_block_stmt_1494/if_stmt_2426__entry__
      -- CP-element group 206: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/$exit
      -- CP-element group 206: 	 branch_block_stmt_1494/if_stmt_2426_dead_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_1494/if_stmt_2426_eval_test/$entry
      -- CP-element group 206: 	 branch_block_stmt_1494/if_stmt_2426_eval_test/$exit
      -- CP-element group 206: 	 branch_block_stmt_1494/if_stmt_2426_eval_test/branch_req
      -- CP-element group 206: 	 branch_block_stmt_1494/R_exitcond_2427_place
      -- CP-element group 206: 	 branch_block_stmt_1494/if_stmt_2426_if_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_1494/if_stmt_2426_else_link/$entry
      -- 
    branch_req_5470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(206), ack => if_stmt_2426_branch_req_0); -- 
    convolution3D_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(167) & convolution3D_CP_3789_elements(205);
      gj_convolution3D_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	349 
    -- CP-element group 207: 	350 
    -- CP-element group 207:  members (24) 
      -- CP-element group 207: 	 branch_block_stmt_1494/merge_stmt_2432__exit__
      -- CP-element group 207: 	 branch_block_stmt_1494/assign_stmt_2439_to_assign_stmt_2454__entry__
      -- CP-element group 207: 	 branch_block_stmt_1494/assign_stmt_2439_to_assign_stmt_2454__exit__
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 207: 	 branch_block_stmt_1494/if_stmt_2426_if_link/$exit
      -- CP-element group 207: 	 branch_block_stmt_1494/if_stmt_2426_if_link/if_choice_transition
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 207: 	 branch_block_stmt_1494/assign_stmt_2439_to_assign_stmt_2454/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/assign_stmt_2439_to_assign_stmt_2454/$exit
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_1494/merge_stmt_2432_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_1494/merge_stmt_2432_PhiAck/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/merge_stmt_2432_PhiAck/$exit
      -- CP-element group 207: 	 branch_block_stmt_1494/merge_stmt_2432_PhiAck/dummy
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2426_branch_ack_1, ack => convolution3D_CP_3789_elements(207)); -- 
    rr_6527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(207), ack => type_cast_2460_inst_req_0); -- 
    cr_6532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(207), ack => type_cast_2460_inst_req_1); -- 
    -- CP-element group 208:  fork  transition  place  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	344 
    -- CP-element group 208: 	345 
    -- CP-element group 208:  members (12) 
      -- CP-element group 208: 	 branch_block_stmt_1494/if_stmt_2426_else_link/$exit
      -- CP-element group 208: 	 branch_block_stmt_1494/if_stmt_2426_else_link/else_choice_transition
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/$entry
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/$entry
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/$entry
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/$entry
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2426_branch_ack_0, ack => convolution3D_CP_3789_elements(208)); -- 
    rr_6484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(208), ack => type_cast_2269_inst_req_0); -- 
    cr_6489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(208), ack => type_cast_2269_inst_req_1); -- 
    -- CP-element group 209:  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	354 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	373 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_1494/if_stmt_2477_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_1494/if_stmt_2477_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_1494/forx_xend215_ifx_xend227
      -- CP-element group 209: 	 branch_block_stmt_1494/forx_xend215_ifx_xend227_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_1494/forx_xend215_ifx_xend227_PhiReq/$exit
      -- 
    if_choice_transition_5500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2477_branch_ack_1, ack => convolution3D_CP_3789_elements(209)); -- 
    -- CP-element group 210:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	354 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (18) 
      -- CP-element group 210: 	 branch_block_stmt_1494/merge_stmt_2483__exit__
      -- CP-element group 210: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499__entry__
      -- CP-element group 210: 	 branch_block_stmt_1494/if_stmt_2477_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_1494/if_stmt_2477_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_1494/forx_xend215_bbx_xnphx_xi356
      -- CP-element group 210: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/$entry
      -- CP-element group 210: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_update_start_
      -- CP-element group 210: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_Update/cr
      -- CP-element group 210: 	 branch_block_stmt_1494/forx_xend215_bbx_xnphx_xi356_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_1494/forx_xend215_bbx_xnphx_xi356_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_1494/merge_stmt_2483_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_1494/merge_stmt_2483_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_1494/merge_stmt_2483_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_1494/merge_stmt_2483_PhiAck/dummy
      -- 
    else_choice_transition_5504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2477_branch_ack_0, ack => convolution3D_CP_3789_elements(210)); -- 
    rr_5517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(210), ack => type_cast_2492_inst_req_0); -- 
    cr_5522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(210), ack => type_cast_2492_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_Sample/ra
      -- 
    ra_5518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2492_inst_ack_0, ack => convolution3D_CP_3789_elements(211)); -- 
    -- CP-element group 212:  fork  transition  place  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	355 
    -- CP-element group 212: 	356 
    -- CP-element group 212:  members (11) 
      -- CP-element group 212: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499__exit__
      -- CP-element group 212: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365
      -- CP-element group 212: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/$exit
      -- CP-element group 212: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_1494/assign_stmt_2489_to_assign_stmt_2499/type_cast_2492_Update/ca
      -- CP-element group 212: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/$entry
      -- CP-element group 212: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/$entry
      -- CP-element group 212: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$entry
      -- 
    ca_5523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2492_inst_ack_1, ack => convolution3D_CP_3789_elements(212)); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	368 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_update_start_
      -- CP-element group 213: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_Sample/ra
      -- CP-element group 213: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_Update/cr
      -- 
    ra_5535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2530_inst_ack_0, ack => convolution3D_CP_3789_elements(213)); -- 
    cr_5539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(213), ack => RPIPE_maxpool_input_pipe_2530_inst_req_1); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_Update/ca
      -- CP-element group 214: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_Sample/rr
      -- 
    ca_5540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2530_inst_ack_1, ack => convolution3D_CP_3789_elements(214)); -- 
    rr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(214), ack => type_cast_2534_inst_req_0); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_Sample/ra
      -- 
    ra_5549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2534_inst_ack_0, ack => convolution3D_CP_3789_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	368 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	219 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_Update/ca
      -- 
    ca_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2534_inst_ack_1, ack => convolution3D_CP_3789_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	368 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_sample_completed_
      -- 
    ra_5563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2549_inst_ack_0, ack => convolution3D_CP_3789_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	368 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_Update/$exit
      -- 
    ca_5568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2549_inst_ack_1, ack => convolution3D_CP_3789_elements(218)); -- 
    -- CP-element group 219:  branch  join  transition  place  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	216 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (10) 
      -- CP-element group 219: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555__exit__
      -- CP-element group 219: 	 branch_block_stmt_1494/if_stmt_2556__entry__
      -- CP-element group 219: 	 branch_block_stmt_1494/if_stmt_2556_eval_test/branch_req
      -- CP-element group 219: 	 branch_block_stmt_1494/if_stmt_2556_eval_test/$exit
      -- CP-element group 219: 	 branch_block_stmt_1494/if_stmt_2556_if_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_1494/if_stmt_2556_eval_test/$entry
      -- CP-element group 219: 	 branch_block_stmt_1494/if_stmt_2556_else_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_1494/if_stmt_2556_dead_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_1494/R_cmpx_xi364_2557_place
      -- CP-element group 219: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/$exit
      -- 
    branch_req_5576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(219), ack => if_stmt_2556_branch_req_0); -- 
    convolution3D_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(216) & convolution3D_CP_3789_elements(218);
      gj_convolution3D_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  place  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	358 
    -- CP-element group 220: 	359 
    -- CP-element group 220: 	361 
    -- CP-element group 220: 	362 
    -- CP-element group 220:  members (20) 
      -- CP-element group 220: 	 branch_block_stmt_1494/if_stmt_2556_if_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365
      -- CP-element group 220: 	 branch_block_stmt_1494/if_stmt_2556_if_link/if_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/Update/cr
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2556_branch_ack_1, ack => convolution3D_CP_3789_elements(220)); -- 
    rr_6600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(220), ack => type_cast_2508_inst_req_0); -- 
    cr_6605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(220), ack => type_cast_2508_inst_req_1); -- 
    rr_6623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(220), ack => type_cast_2515_inst_req_0); -- 
    cr_6628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(220), ack => type_cast_2515_inst_req_1); -- 
    -- CP-element group 221:  fork  transition  place  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	369 
    -- CP-element group 221: 	370 
    -- CP-element group 221:  members (12) 
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373
      -- CP-element group 221: 	 branch_block_stmt_1494/if_stmt_2556_else_link/else_choice_transition
      -- CP-element group 221: 	 branch_block_stmt_1494/if_stmt_2556_else_link/$exit
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/$entry
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/$entry
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/$entry
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/rr
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2556_branch_ack_0, ack => convolution3D_CP_3789_elements(221)); -- 
    rr_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(221), ack => type_cast_2566_inst_req_0); -- 
    cr_6664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(221), ack => type_cast_2566_inst_req_1); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	372 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_Sample/ack
      -- CP-element group 222: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_sample_complete
      -- 
    ack_5616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2595_index_offset_ack_0, ack => convolution3D_CP_3789_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	372 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_request/req
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_Update/$exit
      -- 
    ack_5621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2595_index_offset_ack_1, ack => convolution3D_CP_3789_elements(223)); -- 
    req_5630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(223), ack => addr_of_2596_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_request/ack
      -- CP-element group 224: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_request/$exit
      -- 
    ack_5631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2596_final_reg_ack_0, ack => convolution3D_CP_3789_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	372 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/ptr_deref_2599_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/ptr_deref_2599_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/ptr_deref_2599_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/ptr_deref_2599_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/word_access_start/word_0/rr
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_complete/$exit
      -- 
    ack_5636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2596_final_reg_ack_1, ack => convolution3D_CP_3789_elements(225)); -- 
    rr_5674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(225), ack => ptr_deref_2599_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Sample/word_access_start/word_0/ra
      -- CP-element group 226: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_sample_completed_
      -- 
    ra_5675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2599_store_0_ack_0, ack => convolution3D_CP_3789_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	372 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Update/word_access_complete/word_0/ca
      -- CP-element group 227: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Update/word_access_complete/$exit
      -- 
    ca_5686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2599_store_0_ack_1, ack => convolution3D_CP_3789_elements(227)); -- 
    -- CP-element group 228:  join  transition  place  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	373 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601__exit__
      -- CP-element group 228: 	 branch_block_stmt_1494/getRemainingElementsx_xexit373_ifx_xend227
      -- CP-element group 228: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/$exit
      -- CP-element group 228: 	 branch_block_stmt_1494/getRemainingElementsx_xexit373_ifx_xend227_PhiReq/$entry
      -- CP-element group 228: 	 branch_block_stmt_1494/getRemainingElementsx_xexit373_ifx_xend227_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(222) & convolution3D_CP_3789_elements(227);
      gj_convolution3D_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	373 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_Sample/cra
      -- CP-element group 229: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_sample_completed_
      -- 
    cra_5698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2606_call_ack_0, ack => convolution3D_CP_3789_elements(229)); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	373 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	237 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_Update/cca
      -- CP-element group 230: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_Update/$exit
      -- 
    cca_5703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2606_call_ack_1, ack => convolution3D_CP_3789_elements(230)); -- 
    -- CP-element group 231:  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	373 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (6) 
      -- CP-element group 231: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_Update/req
      -- CP-element group 231: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_Sample/ack
      -- CP-element group 231: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_update_start_
      -- CP-element group 231: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_sample_completed_
      -- 
    ack_5712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2607_inst_ack_0, ack => convolution3D_CP_3789_elements(231)); -- 
    req_5716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(231), ack => WPIPE_output_pipe_2607_inst_req_1); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_Update/ack
      -- CP-element group 232: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_update_completed_
      -- 
    ack_5717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2607_inst_ack_1, ack => convolution3D_CP_3789_elements(232)); -- 
    req_5725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(232), ack => WPIPE_output_pipe_2610_inst_req_0); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_Update/req
      -- CP-element group 233: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_Sample/ack
      -- CP-element group 233: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_update_start_
      -- CP-element group 233: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_sample_completed_
      -- 
    ack_5726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2610_inst_ack_0, ack => convolution3D_CP_3789_elements(233)); -- 
    req_5730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(233), ack => WPIPE_output_pipe_2610_inst_req_1); -- 
    -- CP-element group 234:  transition  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_Update/ack
      -- CP-element group 234: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2610_update_completed_
      -- 
    ack_5731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2610_inst_ack_1, ack => convolution3D_CP_3789_elements(234)); -- 
    req_5739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(234), ack => WPIPE_output_pipe_2613_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_Update/req
      -- CP-element group 235: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_update_start_
      -- CP-element group 235: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_sample_completed_
      -- 
    ack_5740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2613_inst_ack_0, ack => convolution3D_CP_3789_elements(235)); -- 
    req_5744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(235), ack => WPIPE_output_pipe_2613_inst_req_1); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2613_update_completed_
      -- 
    ack_5745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2613_inst_ack_1, ack => convolution3D_CP_3789_elements(236)); -- 
    -- CP-element group 237:  join  fork  transition  place  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: 	230 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237: 	239 
    -- CP-element group 237: 	240 
    -- CP-element group 237: 	241 
    -- CP-element group 237:  members (16) 
      -- CP-element group 237: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615__exit__
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646__entry__
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_Sample/rr
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_Update/cr
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_update_start_
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_update_start_
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/$entry
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_Update/cr
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_Sample/rr
      -- CP-element group 237: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/$exit
      -- 
    rr_5756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(237), ack => type_cast_2630_inst_req_0); -- 
    cr_5761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(237), ack => type_cast_2630_inst_req_1); -- 
    cr_5775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(237), ack => type_cast_2640_inst_req_1); -- 
    rr_5770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(237), ack => type_cast_2640_inst_req_0); -- 
    convolution3D_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(236) & convolution3D_CP_3789_elements(230);
      gj_convolution3D_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_Sample/ra
      -- CP-element group 238: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_sample_completed_
      -- 
    ra_5757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2630_inst_ack_0, ack => convolution3D_CP_3789_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	242 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_Update/ca
      -- CP-element group 239: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2630_update_completed_
      -- 
    ca_5762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2630_inst_ack_1, ack => convolution3D_CP_3789_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	237 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_Sample/ra
      -- CP-element group 240: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_Sample/$exit
      -- 
    ra_5771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2640_inst_ack_0, ack => convolution3D_CP_3789_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	237 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_Update/ca
      -- CP-element group 241: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/type_cast_2640_Update/$exit
      -- 
    ca_5776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2640_inst_ack_1, ack => convolution3D_CP_3789_elements(241)); -- 
    -- CP-element group 242:  join  transition  place  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	239 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	374 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646__exit__
      -- CP-element group 242: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody
      -- CP-element group 242: 	 branch_block_stmt_1494/assign_stmt_2622_to_assign_stmt_2646/$exit
      -- CP-element group 242: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/$entry
      -- CP-element group 242: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2649/$entry
      -- CP-element group 242: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(239) & convolution3D_CP_3789_elements(241);
      gj_convolution3D_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	379 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_Update/req
      -- CP-element group 243: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_update_start_
      -- CP-element group 243: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_sample_completed_
      -- 
    ack_5788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2662_inst_ack_0, ack => convolution3D_CP_3789_elements(243)); -- 
    req_5792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(243), ack => WPIPE_num_out_pipe_2662_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_update_completed_
      -- 
    ack_5793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2662_inst_ack_1, ack => convolution3D_CP_3789_elements(244)); -- 
    req_5801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(244), ack => WPIPE_num_out_pipe_2665_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_Update/req
      -- CP-element group 245: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_update_start_
      -- CP-element group 245: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_sample_completed_
      -- 
    ack_5802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2665_inst_ack_0, ack => convolution3D_CP_3789_elements(245)); -- 
    req_5806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(245), ack => WPIPE_num_out_pipe_2665_inst_req_1); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	251 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2665_update_completed_
      -- 
    ack_5807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2665_inst_ack_1, ack => convolution3D_CP_3789_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	379 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_Sample/cra
      -- CP-element group 247: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_Sample/$exit
      -- 
    cra_5816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2676_call_ack_0, ack => convolution3D_CP_3789_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	379 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	251 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_Update/cca
      -- 
    cca_5821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2676_call_ack_1, ack => convolution3D_CP_3789_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	379 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_Sample/cra
      -- CP-element group 249: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_sample_completed_
      -- 
    cra_5830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2680_call_ack_0, ack => convolution3D_CP_3789_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	379 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_Update/cca
      -- CP-element group 250: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_update_completed_
      -- 
    cca_5835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2680_call_ack_1, ack => convolution3D_CP_3789_elements(250)); -- 
    -- CP-element group 251:  branch  join  transition  place  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	246 
    -- CP-element group 251: 	248 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (10) 
      -- CP-element group 251: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691__exit__
      -- CP-element group 251: 	 branch_block_stmt_1494/if_stmt_2692__entry__
      -- CP-element group 251: 	 branch_block_stmt_1494/R_exitcond5_2693_place
      -- CP-element group 251: 	 branch_block_stmt_1494/if_stmt_2692_else_link/$entry
      -- CP-element group 251: 	 branch_block_stmt_1494/if_stmt_2692_if_link/$entry
      -- CP-element group 251: 	 branch_block_stmt_1494/if_stmt_2692_eval_test/branch_req
      -- CP-element group 251: 	 branch_block_stmt_1494/if_stmt_2692_eval_test/$exit
      -- CP-element group 251: 	 branch_block_stmt_1494/if_stmt_2692_eval_test/$entry
      -- CP-element group 251: 	 branch_block_stmt_1494/if_stmt_2692_dead_link/$entry
      -- CP-element group 251: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/$exit
      -- 
    branch_req_5843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(251), ack => if_stmt_2692_branch_req_0); -- 
    convolution3D_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(246) & convolution3D_CP_3789_elements(248) & convolution3D_CP_3789_elements(250);
      gj_convolution3D_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: 	255 
    -- CP-element group 252: 	256 
    -- CP-element group 252:  members (21) 
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706__entry__
      -- CP-element group 252: 	 branch_block_stmt_1494/merge_stmt_2698__exit__
      -- CP-element group 252: 	 branch_block_stmt_1494/whilex_xbody_whilex_xend
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_update_start_
      -- CP-element group 252: 	 branch_block_stmt_1494/if_stmt_2692_if_link/if_choice_transition
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_1494/if_stmt_2692_if_link/$exit
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/$entry
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_Sample/rr
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_Sample/rr
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_Update/cr
      -- CP-element group 252: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_Update/$entry
      -- CP-element group 252: 	 branch_block_stmt_1494/merge_stmt_2698_PhiAck/dummy
      -- CP-element group 252: 	 branch_block_stmt_1494/merge_stmt_2698_PhiAck/$exit
      -- CP-element group 252: 	 branch_block_stmt_1494/merge_stmt_2698_PhiAck/$entry
      -- CP-element group 252: 	 branch_block_stmt_1494/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 252: 	 branch_block_stmt_1494/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 252: 	 branch_block_stmt_1494/merge_stmt_2698_PhiReqMerge
      -- 
    if_choice_transition_5848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2692_branch_ack_1, ack => convolution3D_CP_3789_elements(252)); -- 
    rr_5865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(252), ack => type_cast_2702_inst_req_0); -- 
    rr_5879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(252), ack => RPIPE_input_done_pipe_2705_inst_req_0); -- 
    cr_5870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(252), ack => type_cast_2702_inst_req_1); -- 
    -- CP-element group 253:  fork  transition  place  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	375 
    -- CP-element group 253: 	376 
    -- CP-element group 253:  members (12) 
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody
      -- CP-element group 253: 	 branch_block_stmt_1494/if_stmt_2692_else_link/$exit
      -- CP-element group 253: 	 branch_block_stmt_1494/if_stmt_2692_else_link/else_choice_transition
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Sample/rr
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/$entry
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/$entry
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/$entry
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/$entry
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Update/cr
      -- CP-element group 253: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Update/$entry
      -- 
    else_choice_transition_5852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2692_branch_ack_0, ack => convolution3D_CP_3789_elements(253)); -- 
    rr_6712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(253), ack => type_cast_2655_inst_req_0); -- 
    cr_6717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(253), ack => type_cast_2655_inst_req_1); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_Sample/ra
      -- 
    ra_5866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2702_inst_ack_0, ack => convolution3D_CP_3789_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	252 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	258 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_Update/ca
      -- CP-element group 255: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/type_cast_2702_Update/$exit
      -- 
    ca_5871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2702_inst_ack_1, ack => convolution3D_CP_3789_elements(255)); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	252 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_Update/cr
      -- CP-element group 256: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_Sample/ra
      -- CP-element group 256: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_update_start_
      -- CP-element group 256: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_sample_completed_
      -- 
    ra_5880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2705_inst_ack_0, ack => convolution3D_CP_3789_elements(256)); -- 
    cr_5884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(256), ack => RPIPE_input_done_pipe_2705_inst_req_1); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_Update/ca
      -- CP-element group 257: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/RPIPE_input_done_pipe_2705_update_completed_
      -- 
    ca_5885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2705_inst_ack_1, ack => convolution3D_CP_3789_elements(257)); -- 
    -- CP-element group 258:  join  transition  place  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	255 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (7) 
      -- CP-element group 258: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706__exit__
      -- CP-element group 258: 	 branch_block_stmt_1494/assign_stmt_2710__entry__
      -- CP-element group 258: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_Sample/rr
      -- CP-element group 258: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_1494/assign_stmt_2703_to_assign_stmt_2706/$exit
      -- CP-element group 258: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_1494/assign_stmt_2710/$entry
      -- 
    rr_5896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(258), ack => RPIPE_input_done_pipe_2709_inst_req_0); -- 
    convolution3D_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(255) & convolution3D_CP_3789_elements(257);
      gj_convolution3D_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_Update/cr
      -- CP-element group 259: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_Sample/ra
      -- CP-element group 259: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_update_start_
      -- CP-element group 259: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_sample_completed_
      -- 
    ra_5897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2709_inst_ack_0, ack => convolution3D_CP_3789_elements(259)); -- 
    cr_5901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(259), ack => RPIPE_input_done_pipe_2709_inst_req_1); -- 
    -- CP-element group 260:  fork  transition  place  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260: 	262 
    -- CP-element group 260: 	264 
    -- CP-element group 260: 	265 
    -- CP-element group 260: 	266 
    -- CP-element group 260: 	267 
    -- CP-element group 260: 	268 
    -- CP-element group 260: 	271 
    -- CP-element group 260:  members (31) 
      -- CP-element group 260: 	 branch_block_stmt_1494/assign_stmt_2710__exit__
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758__entry__
      -- CP-element group 260: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_Update/ca
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/assign_stmt_2710/RPIPE_input_done_pipe_2709_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_update_start_
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_Update/cr
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_update_start_
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/assign_stmt_2710/$exit
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_Update/cr
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_Update/ccr
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_update_start_
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_Update/ccr
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_Sample/crr
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_update_start_
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_update_start_
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_Update/cr
      -- CP-element group 260: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_sample_start_
      -- 
    ca_5902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2709_inst_ack_1, ack => convolution3D_CP_3789_elements(260)); -- 
    rr_5941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(260), ack => type_cast_2726_inst_req_0); -- 
    cr_5932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(260), ack => type_cast_2717_inst_req_1); -- 
    cr_5960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(260), ack => type_cast_2730_inst_req_1); -- 
    ccr_5974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(260), ack => call_stmt_2758_call_req_1); -- 
    ccr_5918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(260), ack => call_stmt_2713_call_req_1); -- 
    rr_5955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(260), ack => type_cast_2730_inst_req_0); -- 
    crr_5913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(260), ack => call_stmt_2713_call_req_0); -- 
    cr_5946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(260), ack => type_cast_2726_inst_req_1); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_Sample/cra
      -- CP-element group 261: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_sample_completed_
      -- 
    cra_5914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2713_call_ack_0, ack => convolution3D_CP_3789_elements(261)); -- 
    -- CP-element group 262:  transition  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (6) 
      -- CP-element group 262: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_Update/cca
      -- CP-element group 262: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2713_update_completed_
      -- 
    cca_5919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2713_call_ack_1, ack => convolution3D_CP_3789_elements(262)); -- 
    rr_5927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(262), ack => type_cast_2717_inst_req_0); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_Sample/ra
      -- CP-element group 263: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_sample_completed_
      -- 
    ra_5928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2717_inst_ack_0, ack => convolution3D_CP_3789_elements(263)); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	260 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	272 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_Update/ca
      -- CP-element group 264: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2717_update_completed_
      -- 
    ca_5933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2717_inst_ack_1, ack => convolution3D_CP_3789_elements(264)); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	260 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_Sample/ra
      -- CP-element group 265: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_sample_completed_
      -- 
    ra_5942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2726_inst_ack_0, ack => convolution3D_CP_3789_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	260 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	269 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_Update/ca
      -- CP-element group 266: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2726_Update/$exit
      -- 
    ca_5947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2726_inst_ack_1, ack => convolution3D_CP_3789_elements(266)); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	260 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_Sample/ra
      -- CP-element group 267: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_sample_completed_
      -- 
    ra_5956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2730_inst_ack_0, ack => convolution3D_CP_3789_elements(267)); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	260 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/type_cast_2730_update_completed_
      -- 
    ca_5961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2730_inst_ack_1, ack => convolution3D_CP_3789_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	266 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_Sample/crr
      -- CP-element group 269: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_sample_start_
      -- 
    crr_5969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(269), ack => call_stmt_2758_call_req_0); -- 
    convolution3D_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(266) & convolution3D_CP_3789_elements(268);
      gj_convolution3D_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_Sample/cra
      -- CP-element group 270: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_sample_completed_
      -- 
    cra_5970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2758_call_ack_0, ack => convolution3D_CP_3789_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	260 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/call_stmt_2758_Update/cca
      -- 
    cca_5975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2758_call_ack_1, ack => convolution3D_CP_3789_elements(271)); -- 
    -- CP-element group 272:  join  fork  transition  place  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	264 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	284 
    -- CP-element group 272: 	285 
    -- CP-element group 272: 	286 
    -- CP-element group 272: 	287 
    -- CP-element group 272: 	288 
    -- CP-element group 272: 	273 
    -- CP-element group 272: 	274 
    -- CP-element group 272: 	275 
    -- CP-element group 272: 	276 
    -- CP-element group 272: 	277 
    -- CP-element group 272: 	278 
    -- CP-element group 272: 	279 
    -- CP-element group 272: 	280 
    -- CP-element group 272: 	281 
    -- CP-element group 272: 	282 
    -- CP-element group 272: 	283 
    -- CP-element group 272:  members (52) 
      -- CP-element group 272: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758__exit__
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857__entry__
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_1494/call_stmt_2713_to_call_stmt_2758/$exit
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_Update/cr
      -- 
    cr_6019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2782_inst_req_1); -- 
    cr_6033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2792_inst_req_1); -- 
    rr_6014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2782_inst_req_0); -- 
    rr_5986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2762_inst_req_0); -- 
    rr_6028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2792_inst_req_0); -- 
    rr_6000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2772_inst_req_0); -- 
    cr_6005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2772_inst_req_1); -- 
    cr_5991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2762_inst_req_1); -- 
    rr_6042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2802_inst_req_0); -- 
    cr_6047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2802_inst_req_1); -- 
    rr_6056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2812_inst_req_0); -- 
    cr_6061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2812_inst_req_1); -- 
    rr_6070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2822_inst_req_0); -- 
    cr_6075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2822_inst_req_1); -- 
    rr_6084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2832_inst_req_0); -- 
    cr_6089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(272), ack => type_cast_2832_inst_req_1); -- 
    convolution3D_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(264) & convolution3D_CP_3789_elements(271);
      gj_convolution3D_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_Sample/ra
      -- CP-element group 273: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_sample_completed_
      -- 
    ra_5987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2762_inst_ack_0, ack => convolution3D_CP_3789_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	309 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_Update/ca
      -- CP-element group 274: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2762_update_completed_
      -- 
    ca_5992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2762_inst_ack_1, ack => convolution3D_CP_3789_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	272 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_Sample/ra
      -- CP-element group 275: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_sample_completed_
      -- 
    ra_6001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_0, ack => convolution3D_CP_3789_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	272 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	306 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2772_Update/ca
      -- 
    ca_6006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_1, ack => convolution3D_CP_3789_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	272 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_Sample/ra
      -- CP-element group 277: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_sample_completed_
      -- 
    ra_6015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2782_inst_ack_0, ack => convolution3D_CP_3789_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	272 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	303 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_Update/ca
      -- CP-element group 278: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2782_Update/$exit
      -- 
    ca_6020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2782_inst_ack_1, ack => convolution3D_CP_3789_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	272 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_sample_completed_
      -- 
    ra_6029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2792_inst_ack_0, ack => convolution3D_CP_3789_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	272 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	300 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2792_Update/ca
      -- 
    ca_6034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2792_inst_ack_1, ack => convolution3D_CP_3789_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	272 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_Sample/ra
      -- 
    ra_6043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_0, ack => convolution3D_CP_3789_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	272 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	297 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2802_Update/ca
      -- 
    ca_6048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_1, ack => convolution3D_CP_3789_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	272 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_sample_completed_
      -- CP-element group 283: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_Sample/ra
      -- 
    ra_6057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2812_inst_ack_0, ack => convolution3D_CP_3789_elements(283)); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	272 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	294 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_update_completed_
      -- CP-element group 284: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2812_Update/ca
      -- 
    ca_6062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2812_inst_ack_1, ack => convolution3D_CP_3789_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	272 
    -- CP-element group 285: successors 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_Sample/ra
      -- 
    ra_6071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_0, ack => convolution3D_CP_3789_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	272 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	291 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2822_Update/ca
      -- 
    ca_6076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_1, ack => convolution3D_CP_3789_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	272 
    -- CP-element group 287: successors 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_Sample/ra
      -- 
    ra_6085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2832_inst_ack_0, ack => convolution3D_CP_3789_elements(287)); -- 
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	272 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/type_cast_2832_Update/ca
      -- CP-element group 288: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_Sample/req
      -- 
    ca_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2832_inst_ack_1, ack => convolution3D_CP_3789_elements(288)); -- 
    req_6098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(288), ack => WPIPE_maxpool_output_pipe_2834_inst_req_0); -- 
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_sample_completed_
      -- CP-element group 289: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_update_start_
      -- CP-element group 289: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_Update/req
      -- 
    ack_6099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2834_inst_ack_0, ack => convolution3D_CP_3789_elements(289)); -- 
    req_6103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(289), ack => WPIPE_maxpool_output_pipe_2834_inst_req_1); -- 
    -- CP-element group 290:  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2834_Update/ack
      -- 
    ack_6104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2834_inst_ack_1, ack => convolution3D_CP_3789_elements(290)); -- 
    -- CP-element group 291:  join  transition  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	286 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_sample_start_
      -- CP-element group 291: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_Sample/$entry
      -- CP-element group 291: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_Sample/req
      -- 
    req_6112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(291), ack => WPIPE_maxpool_output_pipe_2837_inst_req_0); -- 
    convolution3D_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(286) & convolution3D_CP_3789_elements(290);
      gj_convolution3D_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_update_start_
      -- CP-element group 292: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_Sample/ack
      -- CP-element group 292: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_Update/$entry
      -- CP-element group 292: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_Update/req
      -- 
    ack_6113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2837_inst_ack_0, ack => convolution3D_CP_3789_elements(292)); -- 
    req_6117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(292), ack => WPIPE_maxpool_output_pipe_2837_inst_req_1); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2837_Update/ack
      -- 
    ack_6118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2837_inst_ack_1, ack => convolution3D_CP_3789_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	284 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_Sample/req
      -- 
    req_6126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(294), ack => WPIPE_maxpool_output_pipe_2840_inst_req_0); -- 
    convolution3D_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(284) & convolution3D_CP_3789_elements(293);
      gj_convolution3D_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_update_start_
      -- CP-element group 295: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_Update/req
      -- 
    ack_6127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2840_inst_ack_0, ack => convolution3D_CP_3789_elements(295)); -- 
    req_6131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(295), ack => WPIPE_maxpool_output_pipe_2840_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2840_Update/ack
      -- 
    ack_6132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2840_inst_ack_1, ack => convolution3D_CP_3789_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: 	282 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_Sample/req
      -- 
    req_6140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(297), ack => WPIPE_maxpool_output_pipe_2843_inst_req_0); -- 
    convolution3D_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(296) & convolution3D_CP_3789_elements(282);
      gj_convolution3D_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_sample_completed_
      -- CP-element group 298: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_update_start_
      -- CP-element group 298: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_Sample/$exit
      -- CP-element group 298: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_Sample/ack
      -- CP-element group 298: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_Update/req
      -- 
    ack_6141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2843_inst_ack_0, ack => convolution3D_CP_3789_elements(298)); -- 
    req_6145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(298), ack => WPIPE_maxpool_output_pipe_2843_inst_req_1); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_update_completed_
      -- CP-element group 299: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_Update/$exit
      -- CP-element group 299: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2843_Update/ack
      -- 
    ack_6146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2843_inst_ack_1, ack => convolution3D_CP_3789_elements(299)); -- 
    -- CP-element group 300:  join  transition  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: 	280 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_Sample/req
      -- 
    req_6154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(300), ack => WPIPE_maxpool_output_pipe_2846_inst_req_0); -- 
    convolution3D_cp_element_group_300: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_300"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(299) & convolution3D_CP_3789_elements(280);
      gj_convolution3D_cp_element_group_300 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(300), clk => clk, reset => reset); --
    end block;
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_update_start_
      -- CP-element group 301: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_Update/req
      -- 
    ack_6155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2846_inst_ack_0, ack => convolution3D_CP_3789_elements(301)); -- 
    req_6159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(301), ack => WPIPE_maxpool_output_pipe_2846_inst_req_1); -- 
    -- CP-element group 302:  transition  input  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2846_Update/ack
      -- 
    ack_6160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2846_inst_ack_1, ack => convolution3D_CP_3789_elements(302)); -- 
    -- CP-element group 303:  join  transition  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: 	278 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_Sample/req
      -- 
    req_6168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(303), ack => WPIPE_maxpool_output_pipe_2849_inst_req_0); -- 
    convolution3D_cp_element_group_303: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_303"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(302) & convolution3D_CP_3789_elements(278);
      gj_convolution3D_cp_element_group_303 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(303), clk => clk, reset => reset); --
    end block;
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_sample_completed_
      -- CP-element group 304: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_update_start_
      -- CP-element group 304: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_Sample/$exit
      -- CP-element group 304: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_Sample/ack
      -- CP-element group 304: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_Update/req
      -- 
    ack_6169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2849_inst_ack_0, ack => convolution3D_CP_3789_elements(304)); -- 
    req_6173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(304), ack => WPIPE_maxpool_output_pipe_2849_inst_req_1); -- 
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_update_completed_
      -- CP-element group 305: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_Update/$exit
      -- CP-element group 305: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2849_Update/ack
      -- 
    ack_6174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2849_inst_ack_1, ack => convolution3D_CP_3789_elements(305)); -- 
    -- CP-element group 306:  join  transition  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: 	276 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_Sample/req
      -- 
    req_6182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(306), ack => WPIPE_maxpool_output_pipe_2852_inst_req_0); -- 
    convolution3D_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(305) & convolution3D_CP_3789_elements(276);
      gj_convolution3D_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_update_start_
      -- CP-element group 307: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_Update/req
      -- 
    ack_6183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2852_inst_ack_0, ack => convolution3D_CP_3789_elements(307)); -- 
    req_6187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(307), ack => WPIPE_maxpool_output_pipe_2852_inst_req_1); -- 
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2852_Update/ack
      -- 
    ack_6188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2852_inst_ack_1, ack => convolution3D_CP_3789_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: 	274 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_Sample/req
      -- 
    req_6196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(309), ack => WPIPE_maxpool_output_pipe_2855_inst_req_0); -- 
    convolution3D_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(308) & convolution3D_CP_3789_elements(274);
      gj_convolution3D_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_update_start_
      -- CP-element group 310: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_Sample/ack
      -- CP-element group 310: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_Update/req
      -- 
    ack_6197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2855_inst_ack_0, ack => convolution3D_CP_3789_elements(310)); -- 
    req_6201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(310), ack => WPIPE_maxpool_output_pipe_2855_inst_req_1); -- 
    -- CP-element group 311:  transition  place  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311:  members (16) 
      -- CP-element group 311: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857__exit__
      -- CP-element group 311: 	 branch_block_stmt_1494/return__
      -- CP-element group 311: 	 branch_block_stmt_1494/merge_stmt_2859__exit__
      -- CP-element group 311: 	 $exit
      -- CP-element group 311: 	 branch_block_stmt_1494/$exit
      -- CP-element group 311: 	 branch_block_stmt_1494/branch_block_stmt_1494__exit__
      -- CP-element group 311: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/$exit
      -- CP-element group 311: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_1494/merge_stmt_2859_PhiAck/dummy
      -- CP-element group 311: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_1494/assign_stmt_2763_to_assign_stmt_2857/WPIPE_maxpool_output_pipe_2855_Update/ack
      -- CP-element group 311: 	 branch_block_stmt_1494/merge_stmt_2859_PhiAck/$exit
      -- CP-element group 311: 	 branch_block_stmt_1494/merge_stmt_2859_PhiAck/$entry
      -- CP-element group 311: 	 branch_block_stmt_1494/return___PhiReq/$exit
      -- CP-element group 311: 	 branch_block_stmt_1494/return___PhiReq/$entry
      -- CP-element group 311: 	 branch_block_stmt_1494/merge_stmt_2859_PhiReqMerge
      -- 
    ack_6202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2855_inst_ack_1, ack => convolution3D_CP_3789_elements(311)); -- 
    -- CP-element group 312:  transition  output  delay-element  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	86 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	316 
    -- CP-element group 312:  members (5) 
      -- CP-element group 312: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody_PhiReq/$exit
      -- CP-element group 312: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1802/$exit
      -- CP-element group 312: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/$exit
      -- CP-element group 312: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1806_konst_delay_trans
      -- CP-element group 312: 	 branch_block_stmt_1494/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_req
      -- 
    phi_stmt_1802_req_6225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1802_req_6225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(312), ack => phi_stmt_1802_req_0); -- 
    -- Element group convolution3D_CP_3789_elements(312) is a control-delay.
    cp_element_312_delay: control_delay_element  generic map(name => " 312_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(86), ack => convolution3D_CP_3789_elements(312), clk => clk, reset =>reset);
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	128 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313:  members (2) 
      -- CP-element group 313: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Sample/ra
      -- 
    ra_6245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_0, ack => convolution3D_CP_3789_elements(313)); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	128 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (2) 
      -- CP-element group 314: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Update/ca
      -- 
    ca_6250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_1, ack => convolution3D_CP_3789_elements(314)); -- 
    -- CP-element group 315:  join  transition  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (6) 
      -- CP-element group 315: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 315: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/$exit
      -- CP-element group 315: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/$exit
      -- CP-element group 315: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/$exit
      -- CP-element group 315: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/$exit
      -- CP-element group 315: 	 branch_block_stmt_1494/forx_xbody_forx_xbody_PhiReq/phi_stmt_1802/phi_stmt_1802_req
      -- 
    phi_stmt_1802_req_6251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1802_req_6251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(315), ack => phi_stmt_1802_req_1); -- 
    convolution3D_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(313) & convolution3D_CP_3789_elements(314);
      gj_convolution3D_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  merge  transition  place  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	312 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_1494/merge_stmt_1801_PhiReqMerge
      -- CP-element group 316: 	 branch_block_stmt_1494/merge_stmt_1801_PhiAck/$entry
      -- 
    convolution3D_CP_3789_elements(316) <= OrReduce(convolution3D_CP_3789_elements(312) & convolution3D_CP_3789_elements(315));
    -- CP-element group 317:  fork  transition  place  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	122 
    -- CP-element group 317: 	125 
    -- CP-element group 317: 	88 
    -- CP-element group 317: 	90 
    -- CP-element group 317: 	91 
    -- CP-element group 317: 	94 
    -- CP-element group 317: 	98 
    -- CP-element group 317: 	102 
    -- CP-element group 317: 	87 
    -- CP-element group 317: 	106 
    -- CP-element group 317: 	110 
    -- CP-element group 317: 	114 
    -- CP-element group 317: 	118 
    -- CP-element group 317:  members (56) 
      -- CP-element group 317: 	 branch_block_stmt_1494/merge_stmt_1801__exit__
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964__entry__
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Update/word_access_complete/word_0/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Update/word_access_complete/word_0/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Update/word_access_complete/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/ptr_deref_1951_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1943_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1889_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1907_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1925_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_resized_1
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_scaled_1
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_computed_1
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_resize_1/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_resize_1/$exit
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_resize_1/index_resize_req
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_resize_1/index_resize_ack
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_scale_1/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_scale_1/$exit
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_scale_1/scale_rename_req
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_index_scale_1/scale_rename_ack
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_update_start
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_Sample/req
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/array_obj_ref_1814_final_index_sum_regn_Update/req
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_complete/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/addr_of_1815_complete/req
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/RPIPE_maxpool_input_pipe_1818_Sample/rr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1822_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1835_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1853_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_1494/assign_stmt_1816_to_assign_stmt_1964/type_cast_1871_update_start_
      -- CP-element group 317: 	 branch_block_stmt_1494/merge_stmt_1801_PhiAck/$exit
      -- CP-element group 317: 	 branch_block_stmt_1494/merge_stmt_1801_PhiAck/phi_stmt_1802_ack
      -- 
    phi_stmt_1802_ack_6256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1802_ack_0, ack => convolution3D_CP_3789_elements(317)); -- 
    cr_4791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => ptr_deref_1951_store_0_req_1); -- 
    cr_4741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => type_cast_1943_inst_req_1); -- 
    cr_4657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => type_cast_1889_inst_req_1); -- 
    cr_4629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => type_cast_1871_inst_req_1); -- 
    cr_4685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => type_cast_1907_inst_req_1); -- 
    cr_4713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => type_cast_1925_inst_req_1); -- 
    req_4497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => array_obj_ref_1814_index_offset_req_0); -- 
    req_4502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => array_obj_ref_1814_index_offset_req_1); -- 
    req_4517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => addr_of_1815_final_reg_req_1); -- 
    rr_4526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => RPIPE_maxpool_input_pipe_1818_inst_req_0); -- 
    cr_4545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => type_cast_1822_inst_req_1); -- 
    cr_4573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => type_cast_1835_inst_req_1); -- 
    cr_4601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(317), ack => type_cast_1853_inst_req_1); -- 
    -- CP-element group 318:  transition  output  delay-element  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	76 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	322 
    -- CP-element group 318:  members (5) 
      -- CP-element group 318: 	 branch_block_stmt_1494/entry_forx_xend_PhiReq/$exit
      -- CP-element group 318: 	 branch_block_stmt_1494/entry_forx_xend_PhiReq/phi_stmt_1996/$exit
      -- CP-element group 318: 	 branch_block_stmt_1494/entry_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/$exit
      -- CP-element group 318: 	 branch_block_stmt_1494/entry_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_2002_konst_delay_trans
      -- CP-element group 318: 	 branch_block_stmt_1494/entry_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_req
      -- 
    phi_stmt_1996_req_6279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1996_req_6279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(318), ack => phi_stmt_1996_req_1); -- 
    -- Element group convolution3D_CP_3789_elements(318) is a control-delay.
    cp_element_318_delay: control_delay_element  generic map(name => " 318_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(76), ack => convolution3D_CP_3789_elements(318), clk => clk, reset =>reset);
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	127 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (2) 
      -- CP-element group 319: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/Sample/ra
      -- 
    ra_6299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1999_inst_ack_0, ack => convolution3D_CP_3789_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	127 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (2) 
      -- CP-element group 320: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/Update/ca
      -- 
    ca_6304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1999_inst_ack_1, ack => convolution3D_CP_3789_elements(320)); -- 
    -- CP-element group 321:  join  transition  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 321: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/$exit
      -- CP-element group 321: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/$exit
      -- CP-element group 321: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/$exit
      -- CP-element group 321: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_sources/type_cast_1999/SplitProtocol/$exit
      -- CP-element group 321: 	 branch_block_stmt_1494/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1996/phi_stmt_1996_req
      -- 
    phi_stmt_1996_req_6305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1996_req_6305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(321), ack => phi_stmt_1996_req_0); -- 
    convolution3D_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(319) & convolution3D_CP_3789_elements(320);
      gj_convolution3D_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  merge  transition  place  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	318 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (2) 
      -- CP-element group 322: 	 branch_block_stmt_1494/merge_stmt_1995_PhiReqMerge
      -- CP-element group 322: 	 branch_block_stmt_1494/merge_stmt_1995_PhiAck/$entry
      -- 
    convolution3D_CP_3789_elements(322) <= OrReduce(convolution3D_CP_3789_elements(318) & convolution3D_CP_3789_elements(321));
    -- CP-element group 323:  branch  transition  place  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	130 
    -- CP-element group 323: 	129 
    -- CP-element group 323:  members (15) 
      -- CP-element group 323: 	 branch_block_stmt_1494/merge_stmt_1995__exit__
      -- CP-element group 323: 	 branch_block_stmt_1494/assign_stmt_2009_to_assign_stmt_2015__entry__
      -- CP-element group 323: 	 branch_block_stmt_1494/assign_stmt_2009_to_assign_stmt_2015__exit__
      -- CP-element group 323: 	 branch_block_stmt_1494/if_stmt_2016__entry__
      -- CP-element group 323: 	 branch_block_stmt_1494/assign_stmt_2009_to_assign_stmt_2015/$entry
      -- CP-element group 323: 	 branch_block_stmt_1494/assign_stmt_2009_to_assign_stmt_2015/$exit
      -- CP-element group 323: 	 branch_block_stmt_1494/if_stmt_2016_dead_link/$entry
      -- CP-element group 323: 	 branch_block_stmt_1494/if_stmt_2016_else_link/$entry
      -- CP-element group 323: 	 branch_block_stmt_1494/if_stmt_2016_if_link/$entry
      -- CP-element group 323: 	 branch_block_stmt_1494/if_stmt_2016_eval_test/branch_req
      -- CP-element group 323: 	 branch_block_stmt_1494/if_stmt_2016_eval_test/$exit
      -- CP-element group 323: 	 branch_block_stmt_1494/if_stmt_2016_eval_test/$entry
      -- CP-element group 323: 	 branch_block_stmt_1494/R_tobool_2017_place
      -- CP-element group 323: 	 branch_block_stmt_1494/merge_stmt_1995_PhiAck/$exit
      -- CP-element group 323: 	 branch_block_stmt_1494/merge_stmt_1995_PhiAck/phi_stmt_1996_ack
      -- 
    phi_stmt_1996_ack_6310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1996_ack_0, ack => convolution3D_CP_3789_elements(323)); -- 
    branch_req_4825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(323), ack => if_stmt_2016_branch_req_0); -- 
    -- CP-element group 324:  transition  output  delay-element  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	130 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (4) 
      -- CP-element group 324: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/$exit
      -- CP-element group 324: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/$exit
      -- CP-element group 324: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2041_konst_delay_trans
      -- CP-element group 324: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_req
      -- 
    phi_stmt_2037_req_6333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2037_req_6333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(324), ack => phi_stmt_2037_req_0); -- 
    -- Element group convolution3D_CP_3789_elements(324) is a control-delay.
    cp_element_324_delay: control_delay_element  generic map(name => " 324_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(130), ack => convolution3D_CP_3789_elements(324), clk => clk, reset =>reset);
    -- CP-element group 325:  transition  output  delay-element  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	130 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (4) 
      -- CP-element group 325: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/$exit
      -- CP-element group 325: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/$exit
      -- CP-element group 325: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2048_konst_delay_trans
      -- CP-element group 325: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_req
      -- 
    phi_stmt_2044_req_6341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2044_req_6341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(325), ack => phi_stmt_2044_req_0); -- 
    -- Element group convolution3D_CP_3789_elements(325) is a control-delay.
    cp_element_325_delay: control_delay_element  generic map(name => " 325_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(130), ack => convolution3D_CP_3789_elements(325), clk => clk, reset =>reset);
    -- CP-element group 326:  join  transition  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	334 
    -- CP-element group 326:  members (1) 
      -- CP-element group 326: 	 branch_block_stmt_1494/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(324) & convolution3D_CP_3789_elements(325);
      gj_convolution3D_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	138 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (2) 
      -- CP-element group 327: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/Sample/ra
      -- 
    ra_6361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2043_inst_ack_0, ack => convolution3D_CP_3789_elements(327)); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	138 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (2) 
      -- CP-element group 328: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/Update/ca
      -- 
    ca_6366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2043_inst_ack_1, ack => convolution3D_CP_3789_elements(328)); -- 
    -- CP-element group 329:  join  transition  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	333 
    -- CP-element group 329:  members (5) 
      -- CP-element group 329: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/$exit
      -- CP-element group 329: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/$exit
      -- CP-element group 329: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/$exit
      -- CP-element group 329: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_sources/type_cast_2043/SplitProtocol/$exit
      -- CP-element group 329: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2037/phi_stmt_2037_req
      -- 
    phi_stmt_2037_req_6367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2037_req_6367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(329), ack => phi_stmt_2037_req_1); -- 
    convolution3D_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(327) & convolution3D_CP_3789_elements(328);
      gj_convolution3D_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	138 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (2) 
      -- CP-element group 330: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/Sample/ra
      -- 
    ra_6384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2050_inst_ack_0, ack => convolution3D_CP_3789_elements(330)); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	138 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/Update/ca
      -- 
    ca_6389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2050_inst_ack_1, ack => convolution3D_CP_3789_elements(331)); -- 
    -- CP-element group 332:  join  transition  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (5) 
      -- CP-element group 332: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/$exit
      -- CP-element group 332: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/$exit
      -- CP-element group 332: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/$exit
      -- CP-element group 332: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_sources/type_cast_2050/SplitProtocol/$exit
      -- CP-element group 332: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_2044/phi_stmt_2044_req
      -- 
    phi_stmt_2044_req_6390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2044_req_6390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(332), ack => phi_stmt_2044_req_1); -- 
    convolution3D_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(330) & convolution3D_CP_3789_elements(331);
      gj_convolution3D_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  join  transition  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	329 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (1) 
      -- CP-element group 333: 	 branch_block_stmt_1494/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(329) & convolution3D_CP_3789_elements(332);
      gj_convolution3D_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  merge  fork  transition  place  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	326 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (2) 
      -- CP-element group 334: 	 branch_block_stmt_1494/merge_stmt_2036_PhiReqMerge
      -- CP-element group 334: 	 branch_block_stmt_1494/merge_stmt_2036_PhiAck/$entry
      -- 
    convolution3D_CP_3789_elements(334) <= OrReduce(convolution3D_CP_3789_elements(326) & convolution3D_CP_3789_elements(333));
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (1) 
      -- CP-element group 335: 	 branch_block_stmt_1494/merge_stmt_2036_PhiAck/phi_stmt_2037_ack
      -- 
    phi_stmt_2037_ack_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2037_ack_0, ack => convolution3D_CP_3789_elements(335)); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (1) 
      -- CP-element group 336: 	 branch_block_stmt_1494/merge_stmt_2036_PhiAck/phi_stmt_2044_ack
      -- 
    phi_stmt_2044_ack_6396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2044_ack_0, ack => convolution3D_CP_3789_elements(336)); -- 
    -- CP-element group 337:  join  fork  transition  place  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	131 
    -- CP-element group 337: 	134 
    -- CP-element group 337: 	135 
    -- CP-element group 337: 	136 
    -- CP-element group 337:  members (16) 
      -- CP-element group 337: 	 branch_block_stmt_1494/merge_stmt_2036__exit__
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090__entry__
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_update_start_
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/$entry
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2084_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/type_cast_2069_update_start_
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_1494/assign_stmt_2057_to_assign_stmt_2090/RPIPE_maxpool_input_pipe_2065_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_1494/merge_stmt_2036_PhiAck/$exit
      -- 
    rr_4878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(337), ack => type_cast_2084_inst_req_0); -- 
    cr_4883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(337), ack => type_cast_2084_inst_req_1); -- 
    cr_4869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(337), ack => type_cast_2069_inst_req_1); -- 
    rr_4850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(337), ack => RPIPE_maxpool_input_pipe_2065_inst_req_0); -- 
    convolution3D_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(335) & convolution3D_CP_3789_elements(336);
      gj_convolution3D_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	139 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (2) 
      -- CP-element group 338: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/$exit
      -- CP-element group 338: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Sample/ra
      -- 
    ra_6420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2101_inst_ack_0, ack => convolution3D_CP_3789_elements(338)); -- 
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	139 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (2) 
      -- CP-element group 339: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/$exit
      -- CP-element group 339: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/Update/ca
      -- 
    ca_6425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2101_inst_ack_1, ack => convolution3D_CP_3789_elements(339)); -- 
    -- CP-element group 340:  join  transition  place  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (8) 
      -- CP-element group 340: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 340: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/$exit
      -- CP-element group 340: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/$exit
      -- CP-element group 340: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/$exit
      -- CP-element group 340: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_sources/type_cast_2101/SplitProtocol/$exit
      -- CP-element group 340: 	 branch_block_stmt_1494/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_2098/phi_stmt_2098_req
      -- CP-element group 340: 	 branch_block_stmt_1494/merge_stmt_2097_PhiReqMerge
      -- CP-element group 340: 	 branch_block_stmt_1494/merge_stmt_2097_PhiAck/$entry
      -- 
    phi_stmt_2098_req_6426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2098_req_6426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(340), ack => phi_stmt_2098_req_0); -- 
    convolution3D_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(339) & convolution3D_CP_3789_elements(338);
      gj_convolution3D_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	143 
    -- CP-element group 341: 	145 
    -- CP-element group 341: 	140 
    -- CP-element group 341: 	141 
    -- CP-element group 341:  members (29) 
      -- CP-element group 341: 	 branch_block_stmt_1494/merge_stmt_2097__exit__
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136__entry__
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_scale_1/scale_rename_req
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_Update/req
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_resize_1/index_resize_req
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_scale_1/$exit
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_scaled_1
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_complete/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_complete/req
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_scale_1/scale_rename_ack
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_computed_1
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_scale_1/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_resize_1/index_resize_ack
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Update/word_access_complete/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Update/word_access_complete/word_0/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Update/word_access_complete/word_0/cr
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_resize_1/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_resize_1/$exit
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/ptr_deref_2134_update_start_
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_index_resized_1
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/addr_of_2131_update_start_
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_Sample/req
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_update_start
      -- CP-element group 341: 	 branch_block_stmt_1494/assign_stmt_2108_to_assign_stmt_2136/array_obj_ref_2130_final_index_sum_regn_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_1494/merge_stmt_2097_PhiAck/$exit
      -- CP-element group 341: 	 branch_block_stmt_1494/merge_stmt_2097_PhiAck/phi_stmt_2098_ack
      -- 
    phi_stmt_2098_ack_6431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2098_ack_0, ack => convolution3D_CP_3789_elements(341)); -- 
    req_4936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(341), ack => array_obj_ref_2130_index_offset_req_1); -- 
    req_4951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(341), ack => addr_of_2131_final_reg_req_1); -- 
    cr_5001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(341), ack => ptr_deref_2134_store_0_req_1); -- 
    req_4931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(341), ack => array_obj_ref_2130_index_offset_req_0); -- 
    -- CP-element group 342:  merge  fork  transition  place  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	146 
    -- CP-element group 342: 	129 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	147 
    -- CP-element group 342: 	148 
    -- CP-element group 342: 	149 
    -- CP-element group 342: 	150 
    -- CP-element group 342: 	151 
    -- CP-element group 342: 	152 
    -- CP-element group 342:  members (25) 
      -- CP-element group 342: 	 branch_block_stmt_1494/merge_stmt_2138__exit__
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186__entry__
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/$entry
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_update_start_
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_Sample/rr
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_Update/$entry
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2141_Update/cr
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_update_start_
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_Sample/rr
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_Update/$entry
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2145_Update/cr
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_update_start_
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_Sample/rr
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_Update/$entry
      -- CP-element group 342: 	 branch_block_stmt_1494/assign_stmt_2142_to_assign_stmt_2186/type_cast_2149_Update/cr
      -- CP-element group 342: 	 branch_block_stmt_1494/merge_stmt_2138_PhiReqMerge
      -- CP-element group 342: 	 branch_block_stmt_1494/merge_stmt_2138_PhiAck/$entry
      -- CP-element group 342: 	 branch_block_stmt_1494/merge_stmt_2138_PhiAck/$exit
      -- CP-element group 342: 	 branch_block_stmt_1494/merge_stmt_2138_PhiAck/dummy
      -- 
    rr_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(342), ack => type_cast_2141_inst_req_0); -- 
    cr_5018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(342), ack => type_cast_2141_inst_req_1); -- 
    rr_5027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(342), ack => type_cast_2145_inst_req_0); -- 
    cr_5032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(342), ack => type_cast_2145_inst_req_1); -- 
    rr_5041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(342), ack => type_cast_2149_inst_req_0); -- 
    cr_5046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(342), ack => type_cast_2149_inst_req_1); -- 
    convolution3D_CP_3789_elements(342) <= OrReduce(convolution3D_CP_3789_elements(146) & convolution3D_CP_3789_elements(129));
    -- CP-element group 343:  transition  output  delay-element  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	166 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	347 
    -- CP-element group 343:  members (5) 
      -- CP-element group 343: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- CP-element group 343: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_2263/$exit
      -- CP-element group 343: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/$exit
      -- CP-element group 343: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2267_konst_delay_trans
      -- CP-element group 343: 	 branch_block_stmt_1494/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_req
      -- 
    phi_stmt_2263_req_6465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2263_req_6465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(343), ack => phi_stmt_2263_req_0); -- 
    -- Element group convolution3D_CP_3789_elements(343) is a control-delay.
    cp_element_343_delay: control_delay_element  generic map(name => " 343_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(166), ack => convolution3D_CP_3789_elements(343), clk => clk, reset =>reset);
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	208 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (2) 
      -- CP-element group 344: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/Sample/ra
      -- 
    ra_6485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2269_inst_ack_0, ack => convolution3D_CP_3789_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	208 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (2) 
      -- CP-element group 345: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/Update/ca
      -- 
    ca_6490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2269_inst_ack_1, ack => convolution3D_CP_3789_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- CP-element group 346: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/$exit
      -- CP-element group 346: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/$exit
      -- CP-element group 346: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/$exit
      -- CP-element group 346: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2269/SplitProtocol/$exit
      -- CP-element group 346: 	 branch_block_stmt_1494/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_2263/phi_stmt_2263_req
      -- 
    phi_stmt_2263_req_6491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2263_req_6491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(346), ack => phi_stmt_2263_req_1); -- 
    convolution3D_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(344) & convolution3D_CP_3789_elements(345);
      gj_convolution3D_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  merge  transition  place  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	343 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (2) 
      -- CP-element group 347: 	 branch_block_stmt_1494/merge_stmt_2262_PhiReqMerge
      -- CP-element group 347: 	 branch_block_stmt_1494/merge_stmt_2262_PhiAck/$entry
      -- 
    convolution3D_CP_3789_elements(347) <= OrReduce(convolution3D_CP_3789_elements(343) & convolution3D_CP_3789_elements(346));
    -- CP-element group 348:  fork  transition  place  input  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	167 
    -- CP-element group 348: 	202 
    -- CP-element group 348: 	205 
    -- CP-element group 348: 	168 
    -- CP-element group 348: 	170 
    -- CP-element group 348: 	171 
    -- CP-element group 348: 	174 
    -- CP-element group 348: 	178 
    -- CP-element group 348: 	182 
    -- CP-element group 348: 	186 
    -- CP-element group 348: 	190 
    -- CP-element group 348: 	194 
    -- CP-element group 348: 	198 
    -- CP-element group 348:  members (56) 
      -- CP-element group 348: 	 branch_block_stmt_1494/merge_stmt_2262__exit__
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425__entry__
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_resized_1
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_scaled_1
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_computed_1
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_resize_1/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_resize_1/$exit
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_resize_1/index_resize_req
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_resize_1/index_resize_ack
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_scale_1/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_scale_1/$exit
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_scale_1/scale_rename_req
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_index_scale_1/scale_rename_ack
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_update_start
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_Sample/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_Sample/req
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/array_obj_ref_2275_final_index_sum_regn_Update/req
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_complete/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/addr_of_2276_complete/req
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_sample_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_Sample/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/RPIPE_maxpool_input_pipe_2279_Sample/rr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2283_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2296_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2314_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2332_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2350_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2368_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2386_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/type_cast_2404_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Update/word_access_complete/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Update/word_access_complete/word_0/$entry
      -- CP-element group 348: 	 branch_block_stmt_1494/assign_stmt_2277_to_assign_stmt_2425/ptr_deref_2412_Update/word_access_complete/word_0/cr
      -- CP-element group 348: 	 branch_block_stmt_1494/merge_stmt_2262_PhiAck/$exit
      -- CP-element group 348: 	 branch_block_stmt_1494/merge_stmt_2262_PhiAck/phi_stmt_2263_ack
      -- 
    phi_stmt_2263_ack_6496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2263_ack_0, ack => convolution3D_CP_3789_elements(348)); -- 
    req_5167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => array_obj_ref_2275_index_offset_req_0); -- 
    req_5172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => array_obj_ref_2275_index_offset_req_1); -- 
    req_5187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => addr_of_2276_final_reg_req_1); -- 
    rr_5196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => RPIPE_maxpool_input_pipe_2279_inst_req_0); -- 
    cr_5215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => type_cast_2283_inst_req_1); -- 
    cr_5243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => type_cast_2296_inst_req_1); -- 
    cr_5271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => type_cast_2314_inst_req_1); -- 
    cr_5299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => type_cast_2332_inst_req_1); -- 
    cr_5327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => type_cast_2350_inst_req_1); -- 
    cr_5355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => type_cast_2368_inst_req_1); -- 
    cr_5383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => type_cast_2386_inst_req_1); -- 
    cr_5411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => type_cast_2404_inst_req_1); -- 
    cr_5461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(348), ack => ptr_deref_2412_store_0_req_1); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	207 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (2) 
      -- CP-element group 349: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/Sample/ra
      -- 
    ra_6528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_0, ack => convolution3D_CP_3789_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	207 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (2) 
      -- CP-element group 350: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/Update/ca
      -- 
    ca_6533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_1, ack => convolution3D_CP_3789_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (6) 
      -- CP-element group 351: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- CP-element group 351: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/$exit
      -- CP-element group 351: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/$exit
      -- CP-element group 351: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/$exit
      -- CP-element group 351: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2460/SplitProtocol/$exit
      -- CP-element group 351: 	 branch_block_stmt_1494/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_req
      -- 
    phi_stmt_2457_req_6534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2457_req_6534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(351), ack => phi_stmt_2457_req_0); -- 
    convolution3D_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(349) & convolution3D_CP_3789_elements(350);
      gj_convolution3D_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  output  delay-element  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	155 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (5) 
      -- CP-element group 352: 	 branch_block_stmt_1494/ifx_xend_forx_xend215_PhiReq/$exit
      -- CP-element group 352: 	 branch_block_stmt_1494/ifx_xend_forx_xend215_PhiReq/phi_stmt_2457/$exit
      -- CP-element group 352: 	 branch_block_stmt_1494/ifx_xend_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/$exit
      -- CP-element group 352: 	 branch_block_stmt_1494/ifx_xend_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_sources/type_cast_2463_konst_delay_trans
      -- CP-element group 352: 	 branch_block_stmt_1494/ifx_xend_forx_xend215_PhiReq/phi_stmt_2457/phi_stmt_2457_req
      -- 
    phi_stmt_2457_req_6545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2457_req_6545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(352), ack => phi_stmt_2457_req_1); -- 
    -- Element group convolution3D_CP_3789_elements(352) is a control-delay.
    cp_element_352_delay: control_delay_element  generic map(name => " 352_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(155), ack => convolution3D_CP_3789_elements(352), clk => clk, reset =>reset);
    -- CP-element group 353:  merge  transition  place  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (2) 
      -- CP-element group 353: 	 branch_block_stmt_1494/merge_stmt_2456_PhiReqMerge
      -- CP-element group 353: 	 branch_block_stmt_1494/merge_stmt_2456_PhiAck/$entry
      -- 
    convolution3D_CP_3789_elements(353) <= OrReduce(convolution3D_CP_3789_elements(352) & convolution3D_CP_3789_elements(351));
    -- CP-element group 354:  branch  transition  place  input  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	209 
    -- CP-element group 354: 	210 
    -- CP-element group 354:  members (15) 
      -- CP-element group 354: 	 branch_block_stmt_1494/if_stmt_2477__entry__
      -- CP-element group 354: 	 branch_block_stmt_1494/merge_stmt_2456__exit__
      -- CP-element group 354: 	 branch_block_stmt_1494/assign_stmt_2470_to_assign_stmt_2476__entry__
      -- CP-element group 354: 	 branch_block_stmt_1494/assign_stmt_2470_to_assign_stmt_2476__exit__
      -- CP-element group 354: 	 branch_block_stmt_1494/assign_stmt_2470_to_assign_stmt_2476/$entry
      -- CP-element group 354: 	 branch_block_stmt_1494/assign_stmt_2470_to_assign_stmt_2476/$exit
      -- CP-element group 354: 	 branch_block_stmt_1494/if_stmt_2477_dead_link/$entry
      -- CP-element group 354: 	 branch_block_stmt_1494/if_stmt_2477_eval_test/$entry
      -- CP-element group 354: 	 branch_block_stmt_1494/if_stmt_2477_eval_test/$exit
      -- CP-element group 354: 	 branch_block_stmt_1494/if_stmt_2477_eval_test/branch_req
      -- CP-element group 354: 	 branch_block_stmt_1494/R_tobool218_2478_place
      -- CP-element group 354: 	 branch_block_stmt_1494/if_stmt_2477_if_link/$entry
      -- CP-element group 354: 	 branch_block_stmt_1494/if_stmt_2477_else_link/$entry
      -- CP-element group 354: 	 branch_block_stmt_1494/merge_stmt_2456_PhiAck/$exit
      -- CP-element group 354: 	 branch_block_stmt_1494/merge_stmt_2456_PhiAck/phi_stmt_2457_ack
      -- 
    phi_stmt_2457_ack_6550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2457_ack_0, ack => convolution3D_CP_3789_elements(354)); -- 
    branch_req_5495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(354), ack => if_stmt_2477_branch_req_0); -- 
    -- CP-element group 355:  transition  output  delay-element  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	212 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (4) 
      -- CP-element group 355: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/$exit
      -- CP-element group 355: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/$exit
      -- CP-element group 355: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2506_konst_delay_trans
      -- CP-element group 355: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_req
      -- 
    phi_stmt_2502_req_6573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2502_req_6573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(355), ack => phi_stmt_2502_req_0); -- 
    -- Element group convolution3D_CP_3789_elements(355) is a control-delay.
    cp_element_355_delay: control_delay_element  generic map(name => " 355_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(212), ack => convolution3D_CP_3789_elements(355), clk => clk, reset =>reset);
    -- CP-element group 356:  transition  output  delay-element  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	212 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (4) 
      -- CP-element group 356: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/$exit
      -- CP-element group 356: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$exit
      -- CP-element group 356: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2513_konst_delay_trans
      -- CP-element group 356: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_req
      -- 
    phi_stmt_2509_req_6581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2509_req_6581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(356), ack => phi_stmt_2509_req_0); -- 
    -- Element group convolution3D_CP_3789_elements(356) is a control-delay.
    cp_element_356_delay: control_delay_element  generic map(name => " 356_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(212), ack => convolution3D_CP_3789_elements(356), clk => clk, reset =>reset);
    -- CP-element group 357:  join  transition  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	365 
    -- CP-element group 357:  members (1) 
      -- CP-element group 357: 	 branch_block_stmt_1494/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(355) & convolution3D_CP_3789_elements(356);
      gj_convolution3D_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  transition  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	220 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (2) 
      -- CP-element group 358: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/Sample/ra
      -- 
    ra_6601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_0, ack => convolution3D_CP_3789_elements(358)); -- 
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	220 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (2) 
      -- CP-element group 359: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/Update/ca
      -- 
    ca_6606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_1, ack => convolution3D_CP_3789_elements(359)); -- 
    -- CP-element group 360:  join  transition  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	364 
    -- CP-element group 360:  members (5) 
      -- CP-element group 360: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/$exit
      -- CP-element group 360: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/$exit
      -- CP-element group 360: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/$exit
      -- CP-element group 360: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_sources/type_cast_2508/SplitProtocol/$exit
      -- CP-element group 360: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2502/phi_stmt_2502_req
      -- 
    phi_stmt_2502_req_6607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2502_req_6607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(360), ack => phi_stmt_2502_req_1); -- 
    convolution3D_cp_element_group_360: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_360"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(358) & convolution3D_CP_3789_elements(359);
      gj_convolution3D_cp_element_group_360 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(360), clk => clk, reset => reset); --
    end block;
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	220 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (2) 
      -- CP-element group 361: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/Sample/ra
      -- 
    ra_6624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2515_inst_ack_0, ack => convolution3D_CP_3789_elements(361)); -- 
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	220 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/Update/ca
      -- 
    ca_6629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2515_inst_ack_1, ack => convolution3D_CP_3789_elements(362)); -- 
    -- CP-element group 363:  join  transition  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/$exit
      -- CP-element group 363: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/$exit
      -- CP-element group 363: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/$exit
      -- CP-element group 363: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_sources/type_cast_2515/SplitProtocol/$exit
      -- CP-element group 363: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2509/phi_stmt_2509_req
      -- 
    phi_stmt_2509_req_6630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2509_req_6630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(363), ack => phi_stmt_2509_req_1); -- 
    convolution3D_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(361) & convolution3D_CP_3789_elements(362);
      gj_convolution3D_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  join  transition  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	360 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (1) 
      -- CP-element group 364: 	 branch_block_stmt_1494/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(360) & convolution3D_CP_3789_elements(363);
      gj_convolution3D_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  merge  fork  transition  place  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	357 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: 	367 
    -- CP-element group 365:  members (2) 
      -- CP-element group 365: 	 branch_block_stmt_1494/merge_stmt_2501_PhiReqMerge
      -- CP-element group 365: 	 branch_block_stmt_1494/merge_stmt_2501_PhiAck/$entry
      -- 
    convolution3D_CP_3789_elements(365) <= OrReduce(convolution3D_CP_3789_elements(357) & convolution3D_CP_3789_elements(364));
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (1) 
      -- CP-element group 366: 	 branch_block_stmt_1494/merge_stmt_2501_PhiAck/phi_stmt_2502_ack
      -- 
    phi_stmt_2502_ack_6635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2502_ack_0, ack => convolution3D_CP_3789_elements(366)); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	365 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (1) 
      -- CP-element group 367: 	 branch_block_stmt_1494/merge_stmt_2501_PhiAck/phi_stmt_2509_ack
      -- 
    phi_stmt_2509_ack_6636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2509_ack_0, ack => convolution3D_CP_3789_elements(367)); -- 
    -- CP-element group 368:  join  fork  transition  place  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	213 
    -- CP-element group 368: 	216 
    -- CP-element group 368: 	217 
    -- CP-element group 368: 	218 
    -- CP-element group 368:  members (16) 
      -- CP-element group 368: 	 branch_block_stmt_1494/merge_stmt_2501__exit__
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555__entry__
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_Sample/rr
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_update_start_
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2549_sample_start_
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/$entry
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_sample_start_
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/RPIPE_maxpool_input_pipe_2530_Sample/rr
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_update_start_
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_1494/assign_stmt_2522_to_assign_stmt_2555/type_cast_2534_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_1494/merge_stmt_2501_PhiAck/$exit
      -- 
    rr_5562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(368), ack => type_cast_2549_inst_req_0); -- 
    cr_5567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(368), ack => type_cast_2549_inst_req_1); -- 
    rr_5534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(368), ack => RPIPE_maxpool_input_pipe_2530_inst_req_0); -- 
    cr_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(368), ack => type_cast_2534_inst_req_1); -- 
    convolution3D_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(366) & convolution3D_CP_3789_elements(367);
      gj_convolution3D_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	221 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	371 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/ra
      -- 
    ra_6660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2566_inst_ack_0, ack => convolution3D_CP_3789_elements(369)); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	221 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (2) 
      -- CP-element group 370: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/ca
      -- 
    ca_6665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2566_inst_ack_1, ack => convolution3D_CP_3789_elements(370)); -- 
    -- CP-element group 371:  join  transition  place  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (8) 
      -- CP-element group 371: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/$exit
      -- CP-element group 371: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/$exit
      -- CP-element group 371: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$exit
      -- CP-element group 371: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/$exit
      -- CP-element group 371: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/$exit
      -- CP-element group 371: 	 branch_block_stmt_1494/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2563/phi_stmt_2563_req
      -- CP-element group 371: 	 branch_block_stmt_1494/merge_stmt_2562_PhiReqMerge
      -- CP-element group 371: 	 branch_block_stmt_1494/merge_stmt_2562_PhiAck/$entry
      -- 
    phi_stmt_2563_req_6666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2563_req_6666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(371), ack => phi_stmt_2563_req_0); -- 
    convolution3D_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(369) & convolution3D_CP_3789_elements(370);
      gj_convolution3D_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	222 
    -- CP-element group 372: 	223 
    -- CP-element group 372: 	225 
    -- CP-element group 372: 	227 
    -- CP-element group 372:  members (29) 
      -- CP-element group 372: 	 branch_block_stmt_1494/merge_stmt_2562__exit__
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601__entry__
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_computed_1
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_scale_1/scale_rename_ack
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_resized_1
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_scale_1/$exit
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_scale_1/scale_rename_req
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_scaled_1
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_resize_1/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_resize_1/$exit
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_update_start_
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_update_start_
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_complete/req
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/addr_of_2596_complete/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_Update/req
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_scale_1/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_resize_1/index_resize_ack
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_index_resize_1/index_resize_req
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_Sample/req
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Update/word_access_complete/word_0/cr
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Update/word_access_complete/word_0/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/array_obj_ref_2595_final_index_sum_regn_update_start
      -- CP-element group 372: 	 branch_block_stmt_1494/assign_stmt_2573_to_assign_stmt_2601/ptr_deref_2599_Update/word_access_complete/$entry
      -- CP-element group 372: 	 branch_block_stmt_1494/merge_stmt_2562_PhiAck/$exit
      -- CP-element group 372: 	 branch_block_stmt_1494/merge_stmt_2562_PhiAck/phi_stmt_2563_ack
      -- 
    phi_stmt_2563_ack_6671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2563_ack_0, ack => convolution3D_CP_3789_elements(372)); -- 
    req_5635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(372), ack => addr_of_2596_final_reg_req_1); -- 
    req_5620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(372), ack => array_obj_ref_2595_index_offset_req_1); -- 
    req_5615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(372), ack => array_obj_ref_2595_index_offset_req_0); -- 
    cr_5685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(372), ack => ptr_deref_2599_store_0_req_1); -- 
    -- CP-element group 373:  merge  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	209 
    -- CP-element group 373: 	228 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	229 
    -- CP-element group 373: 	230 
    -- CP-element group 373: 	231 
    -- CP-element group 373:  members (16) 
      -- CP-element group 373: 	 branch_block_stmt_1494/merge_stmt_2603__exit__
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615__entry__
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_Sample/crr
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_update_start_
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_Sample/req
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/WPIPE_output_pipe_2607_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_Update/ccr
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/call_stmt_2606_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_1494/call_stmt_2606_to_assign_stmt_2615/$entry
      -- CP-element group 373: 	 branch_block_stmt_1494/merge_stmt_2603_PhiReqMerge
      -- CP-element group 373: 	 branch_block_stmt_1494/merge_stmt_2603_PhiAck/$entry
      -- CP-element group 373: 	 branch_block_stmt_1494/merge_stmt_2603_PhiAck/$exit
      -- CP-element group 373: 	 branch_block_stmt_1494/merge_stmt_2603_PhiAck/dummy
      -- 
    crr_5697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(373), ack => call_stmt_2606_call_req_0); -- 
    req_5711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(373), ack => WPIPE_output_pipe_2607_inst_req_0); -- 
    ccr_5702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(373), ack => call_stmt_2606_call_req_1); -- 
    convolution3D_CP_3789_elements(373) <= OrReduce(convolution3D_CP_3789_elements(209) & convolution3D_CP_3789_elements(228));
    -- CP-element group 374:  transition  output  delay-element  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	242 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	378 
    -- CP-element group 374:  members (5) 
      -- CP-element group 374: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_req
      -- CP-element group 374: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2653_konst_delay_trans
      -- CP-element group 374: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/$exit
      -- CP-element group 374: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2649/$exit
      -- CP-element group 374: 	 branch_block_stmt_1494/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_2649_req_6693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2649_req_6693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(374), ack => phi_stmt_2649_req_0); -- 
    -- Element group convolution3D_CP_3789_elements(374) is a control-delay.
    cp_element_374_delay: control_delay_element  generic map(name => " 374_delay", delay_value => 1)  port map(req => convolution3D_CP_3789_elements(242), ack => convolution3D_CP_3789_elements(374), clk => clk, reset =>reset);
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	253 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (2) 
      -- CP-element group 375: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Sample/ra
      -- CP-element group 375: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Sample/$exit
      -- 
    ra_6713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_0, ack => convolution3D_CP_3789_elements(375)); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	253 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (2) 
      -- CP-element group 376: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Update/ca
      -- CP-element group 376: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/Update/$exit
      -- 
    ca_6718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_1, ack => convolution3D_CP_3789_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (6) 
      -- CP-element group 377: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/SplitProtocol/$exit
      -- CP-element group 377: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/type_cast_2655/$exit
      -- CP-element group 377: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_sources/$exit
      -- CP-element group 377: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/$exit
      -- CP-element group 377: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 377: 	 branch_block_stmt_1494/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2649/phi_stmt_2649_req
      -- 
    phi_stmt_2649_req_6719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2649_req_6719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(377), ack => phi_stmt_2649_req_1); -- 
    convolution3D_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3789_elements(375) & convolution3D_CP_3789_elements(376);
      gj_convolution3D_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3789_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  merge  transition  place  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	374 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (2) 
      -- CP-element group 378: 	 branch_block_stmt_1494/merge_stmt_2648_PhiAck/$entry
      -- CP-element group 378: 	 branch_block_stmt_1494/merge_stmt_2648_PhiReqMerge
      -- 
    convolution3D_CP_3789_elements(378) <= OrReduce(convolution3D_CP_3789_elements(374) & convolution3D_CP_3789_elements(377));
    -- CP-element group 379:  fork  transition  place  input  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	243 
    -- CP-element group 379: 	247 
    -- CP-element group 379: 	248 
    -- CP-element group 379: 	249 
    -- CP-element group 379: 	250 
    -- CP-element group 379:  members (20) 
      -- CP-element group 379: 	 branch_block_stmt_1494/merge_stmt_2648__exit__
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691__entry__
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_update_start_
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_Sample/crr
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_Update/ccr
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2676_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_Update/ccr
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_Sample/req
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_Sample/crr
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/WPIPE_num_out_pipe_2662_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_update_start_
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/$entry
      -- CP-element group 379: 	 branch_block_stmt_1494/assign_stmt_2661_to_assign_stmt_2691/call_stmt_2680_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_1494/merge_stmt_2648_PhiAck/phi_stmt_2649_ack
      -- CP-element group 379: 	 branch_block_stmt_1494/merge_stmt_2648_PhiAck/$exit
      -- 
    phi_stmt_2649_ack_6724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2649_ack_0, ack => convolution3D_CP_3789_elements(379)); -- 
    crr_5815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(379), ack => call_stmt_2676_call_req_0); -- 
    ccr_5820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(379), ack => call_stmt_2676_call_req_1); -- 
    ccr_5834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(379), ack => call_stmt_2680_call_req_1); -- 
    req_5787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(379), ack => WPIPE_num_out_pipe_2662_inst_req_0); -- 
    crr_5829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3789_elements(379), ack => call_stmt_2680_call_req_0); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1991_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_2178_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_2452_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_2754_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_2108 : std_logic_vector(63 downto 0);
    signal R_indvar411_2274_resized : std_logic_vector(13 downto 0);
    signal R_indvar411_2274_scaled : std_logic_vector(13 downto 0);
    signal R_indvar425_1813_resized : std_logic_vector(13 downto 0);
    signal R_indvar425_1813_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_2129_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_2129_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_2594_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_2594_scaled : std_logic_vector(13 downto 0);
    signal add102_1859 : std_logic_vector(63 downto 0);
    signal add108_1877 : std_logic_vector(63 downto 0);
    signal add114_1895 : std_logic_vector(63 downto 0);
    signal add120_1913 : std_logic_vector(63 downto 0);
    signal add1216x_xi370_2579 : std_logic_vector(63 downto 0);
    signal add1216x_xi_2114 : std_logic_vector(63 downto 0);
    signal add126_1931 : std_logic_vector(63 downto 0);
    signal add132_1949 : std_logic_vector(63 downto 0);
    signal add13_1544 : std_logic_vector(15 downto 0);
    signal add171_2302 : std_logic_vector(63 downto 0);
    signal add177_2320 : std_logic_vector(63 downto 0);
    signal add183_2338 : std_logic_vector(63 downto 0);
    signal add189_2356 : std_logic_vector(63 downto 0);
    signal add195_2374 : std_logic_vector(63 downto 0);
    signal add201_2392 : std_logic_vector(63 downto 0);
    signal add207_2410 : std_logic_vector(63 downto 0);
    signal add23_1569 : std_logic_vector(15 downto 0);
    signal add33_1594 : std_logic_vector(15 downto 0);
    signal add43_1619 : std_logic_vector(15 downto 0);
    signal add53_1644 : std_logic_vector(15 downto 0);
    signal add63_1669 : std_logic_vector(63 downto 0);
    signal add73_1694 : std_logic_vector(15 downto 0);
    signal add96_1841 : std_logic_vector(63 downto 0);
    signal add_1519 : std_logic_vector(31 downto 0);
    signal addx_xi361_2540 : std_logic_vector(63 downto 0);
    signal addx_xi_2075 : std_logic_vector(63 downto 0);
    signal and217_2470 : std_logic_vector(63 downto 0);
    signal and_2009 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1814_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1814_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1814_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1814_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1814_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1814_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2130_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2130_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2130_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2130_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2130_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2130_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2275_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2275_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2275_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2275_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2275_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2275_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2595_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2595_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2595_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2595_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2595_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2595_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_2132 : std_logic_vector(31 downto 0);
    signal arrayidx211_2277 : std_logic_vector(31 downto 0);
    signal arrayidx226_2597 : std_logic_vector(31 downto 0);
    signal arrayidx_1816 : std_logic_vector(31 downto 0);
    signal call105_1868 : std_logic_vector(7 downto 0);
    signal call111_1886 : std_logic_vector(7 downto 0);
    signal call117_1904 : std_logic_vector(7 downto 0);
    signal call11_1535 : std_logic_vector(7 downto 0);
    signal call123_1922 : std_logic_vector(7 downto 0);
    signal call129_1940 : std_logic_vector(7 downto 0);
    signal call164_2280 : std_logic_vector(7 downto 0);
    signal call168_2293 : std_logic_vector(7 downto 0);
    signal call16_1547 : std_logic_vector(7 downto 0);
    signal call174_2311 : std_logic_vector(7 downto 0);
    signal call180_2329 : std_logic_vector(7 downto 0);
    signal call186_2347 : std_logic_vector(7 downto 0);
    signal call192_2365 : std_logic_vector(7 downto 0);
    signal call198_2383 : std_logic_vector(7 downto 0);
    signal call204_2401 : std_logic_vector(7 downto 0);
    signal call21_1560 : std_logic_vector(7 downto 0);
    signal call229_2606 : std_logic_vector(63 downto 0);
    signal call26_1572 : std_logic_vector(7 downto 0);
    signal call270_2706 : std_logic_vector(7 downto 0);
    signal call273_2710 : std_logic_vector(7 downto 0);
    signal call275_2713 : std_logic_vector(63 downto 0);
    signal call2_1510 : std_logic_vector(7 downto 0);
    signal call31_1585 : std_logic_vector(7 downto 0);
    signal call36_1597 : std_logic_vector(7 downto 0);
    signal call41_1610 : std_logic_vector(7 downto 0);
    signal call46_1622 : std_logic_vector(7 downto 0);
    signal call51_1635 : std_logic_vector(7 downto 0);
    signal call56_1647 : std_logic_vector(7 downto 0);
    signal call61_1660 : std_logic_vector(7 downto 0);
    signal call66_1672 : std_logic_vector(7 downto 0);
    signal call6_1522 : std_logic_vector(7 downto 0);
    signal call71_1685 : std_logic_vector(7 downto 0);
    signal call89_1819 : std_logic_vector(7 downto 0);
    signal call93_1832 : std_logic_vector(7 downto 0);
    signal call99_1850 : std_logic_vector(7 downto 0);
    signal call_1497 : std_logic_vector(7 downto 0);
    signal callx_xi359_2531 : std_logic_vector(7 downto 0);
    signal callx_xi_2066 : std_logic_vector(7 downto 0);
    signal cmp161379_2186 : std_logic_vector(0 downto 0);
    signal cmp383_1723 : std_logic_vector(0 downto 0);
    signal cmpx_xi364_2555 : std_logic_vector(0 downto 0);
    signal cmpx_xi_2090 : std_logic_vector(0 downto 0);
    signal conv101_1854 : std_logic_vector(63 downto 0);
    signal conv107_1872 : std_logic_vector(63 downto 0);
    signal conv113_1890 : std_logic_vector(63 downto 0);
    signal conv119_1908 : std_logic_vector(63 downto 0);
    signal conv125_1926 : std_logic_vector(63 downto 0);
    signal conv12_1539 : std_logic_vector(15 downto 0);
    signal conv131_1944 : std_logic_vector(63 downto 0);
    signal conv145_2142 : std_logic_vector(63 downto 0);
    signal conv147_2146 : std_logic_vector(63 downto 0);
    signal conv153_2150 : std_logic_vector(63 downto 0);
    signal conv155_2180 : std_logic_vector(63 downto 0);
    signal conv165_2284 : std_logic_vector(63 downto 0);
    signal conv170_2297 : std_logic_vector(63 downto 0);
    signal conv176_2315 : std_logic_vector(63 downto 0);
    signal conv182_2333 : std_logic_vector(63 downto 0);
    signal conv188_2351 : std_logic_vector(63 downto 0);
    signal conv194_2369 : std_logic_vector(63 downto 0);
    signal conv19_1551 : std_logic_vector(15 downto 0);
    signal conv1_1501 : std_logic_vector(31 downto 0);
    signal conv200_2387 : std_logic_vector(63 downto 0);
    signal conv206_2405 : std_logic_vector(63 downto 0);
    signal conv22_1564 : std_logic_vector(15 downto 0);
    signal conv230_2703 : std_logic_vector(63 downto 0);
    signal conv254_2673 : std_logic_vector(63 downto 0);
    signal conv276_2718 : std_logic_vector(63 downto 0);
    signal conv281_2727 : std_logic_vector(63 downto 0);
    signal conv283_2731 : std_logic_vector(63 downto 0);
    signal conv288_2756 : std_logic_vector(63 downto 0);
    signal conv292_2763 : std_logic_vector(7 downto 0);
    signal conv298_2773 : std_logic_vector(7 downto 0);
    signal conv29_1576 : std_logic_vector(15 downto 0);
    signal conv2x_xi354_2493 : std_logic_vector(31 downto 0);
    signal conv2x_xi_2028 : std_logic_vector(31 downto 0);
    signal conv304_2783 : std_logic_vector(7 downto 0);
    signal conv310_2793 : std_logic_vector(7 downto 0);
    signal conv316_2803 : std_logic_vector(7 downto 0);
    signal conv322_2813 : std_logic_vector(7 downto 0);
    signal conv328_2823 : std_logic_vector(7 downto 0);
    signal conv32_1589 : std_logic_vector(15 downto 0);
    signal conv334_2833 : std_logic_vector(7 downto 0);
    signal conv39_1601 : std_logic_vector(15 downto 0);
    signal conv3_1514 : std_logic_vector(31 downto 0);
    signal conv42_1614 : std_logic_vector(15 downto 0);
    signal conv49_1626 : std_logic_vector(15 downto 0);
    signal conv52_1639 : std_logic_vector(15 downto 0);
    signal conv59_1651 : std_logic_vector(63 downto 0);
    signal conv5x_xi360_2535 : std_logic_vector(63 downto 0);
    signal conv5x_xi_2070 : std_logic_vector(63 downto 0);
    signal conv62_1664 : std_logic_vector(63 downto 0);
    signal conv69_1676 : std_logic_vector(15 downto 0);
    signal conv72_1689 : std_logic_vector(15 downto 0);
    signal conv79_1698 : std_logic_vector(31 downto 0);
    signal conv81_1702 : std_logic_vector(31 downto 0);
    signal conv83_1717 : std_logic_vector(63 downto 0);
    signal conv90_1823 : std_logic_vector(63 downto 0);
    signal conv95_1836 : std_logic_vector(63 downto 0);
    signal conv9_1526 : std_logic_vector(15 downto 0);
    signal convx_xi363_2550 : std_logic_vector(31 downto 0);
    signal convx_xi_2085 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi358_2509 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_2044 : std_logic_vector(63 downto 0);
    signal exitcond28_1964 : std_logic_vector(0 downto 0);
    signal exitcond5_2691 : std_logic_vector(0 downto 0);
    signal exitcond_2425 : std_logic_vector(0 downto 0);
    signal iNsTr_34_2063 : std_logic_vector(15 downto 0);
    signal iNsTr_56_2489 : std_logic_vector(63 downto 0);
    signal iNsTr_68_2528 : std_logic_vector(15 downto 0);
    signal iNsTr_94_2573 : std_logic_vector(63 downto 0);
    signal indvar411_2263 : std_logic_vector(63 downto 0);
    signal indvar425_1802 : std_logic_vector(63 downto 0);
    signal indvar_2649 : std_logic_vector(63 downto 0);
    signal indvarx_xnext412_2420 : std_logic_vector(63 downto 0);
    signal indvarx_xnext426_1959 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_2686 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_1996 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_2457 : std_logic_vector(63 downto 0);
    signal mul148_2155 : std_logic_vector(63 downto 0);
    signal mul151_2160 : std_logic_vector(63 downto 0);
    signal mul154_2165 : std_logic_vector(63 downto 0);
    signal mul253_2661 : std_logic_vector(63 downto 0);
    signal mul284_2737 : std_logic_vector(63 downto 0);
    signal mul287_2742 : std_logic_vector(63 downto 0);
    signal mul82_1712 : std_logic_vector(31 downto 0);
    signal mul_1707 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi357_2502 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_2037 : std_logic_vector(15 downto 0);
    signal phitmp387_2454 : std_logic_vector(63 downto 0);
    signal phitmp_1993 : std_logic_vector(63 downto 0);
    signal ptr_deref_1951_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1951_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1951_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1951_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1951_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1951_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2134_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2134_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2134_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2134_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2134_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2134_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2412_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2412_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2412_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2412_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2412_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2412_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2599_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2599_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2599_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2599_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2599_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2599_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext352_2747 : std_logic_vector(63 downto 0);
    signal sext_2171 : std_logic_vector(63 downto 0);
    signal sh_promx_xi371_2585 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_2120 : std_logic_vector(63 downto 0);
    signal shl104_1865 : std_logic_vector(63 downto 0);
    signal shl10_1532 : std_logic_vector(15 downto 0);
    signal shl110_1883 : std_logic_vector(63 downto 0);
    signal shl116_1901 : std_logic_vector(63 downto 0);
    signal shl122_1919 : std_logic_vector(63 downto 0);
    signal shl128_1937 : std_logic_vector(63 downto 0);
    signal shl14x_xi372_2590 : std_logic_vector(63 downto 0);
    signal shl14x_xi_2125 : std_logic_vector(63 downto 0);
    signal shl167_2290 : std_logic_vector(63 downto 0);
    signal shl173_2308 : std_logic_vector(63 downto 0);
    signal shl179_2326 : std_logic_vector(63 downto 0);
    signal shl185_2344 : std_logic_vector(63 downto 0);
    signal shl191_2362 : std_logic_vector(63 downto 0);
    signal shl197_2380 : std_logic_vector(63 downto 0);
    signal shl203_2398 : std_logic_vector(63 downto 0);
    signal shl20_1557 : std_logic_vector(15 downto 0);
    signal shl30_1582 : std_logic_vector(15 downto 0);
    signal shl40_1607 : std_logic_vector(15 downto 0);
    signal shl50_1632 : std_logic_vector(15 downto 0);
    signal shl60_1657 : std_logic_vector(63 downto 0);
    signal shl70_1682 : std_logic_vector(15 downto 0);
    signal shl8x_xi362_2546 : std_logic_vector(63 downto 0);
    signal shl8x_xi362x_xlcssa_2563 : std_logic_vector(63 downto 0);
    signal shl8x_xi_2081 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_2098 : std_logic_vector(63 downto 0);
    signal shl92_1829 : std_logic_vector(63 downto 0);
    signal shl98_1847 : std_logic_vector(63 downto 0);
    signal shl_1507 : std_logic_vector(31 downto 0);
    signal shlx_xi355_2499 : std_logic_vector(31 downto 0);
    signal shlx_xi_2034 : std_logic_vector(31 downto 0);
    signal shr295_2769 : std_logic_vector(63 downto 0);
    signal shr301_2779 : std_logic_vector(63 downto 0);
    signal shr307_2789 : std_logic_vector(63 downto 0);
    signal shr313_2799 : std_logic_vector(63 downto 0);
    signal shr319_2809 : std_logic_vector(63 downto 0);
    signal shr325_2819 : std_logic_vector(63 downto 0);
    signal shr331_2829 : std_logic_vector(63 downto 0);
    signal sub_2723 : std_logic_vector(63 downto 0);
    signal tmp10_2214 : std_logic_vector(63 downto 0);
    signal tmp11_2218 : std_logic_vector(63 downto 0);
    signal tmp12_2223 : std_logic_vector(63 downto 0);
    signal tmp13_2227 : std_logic_vector(63 downto 0);
    signal tmp14_2232 : std_logic_vector(63 downto 0);
    signal tmp15_2236 : std_logic_vector(31 downto 0);
    signal tmp16_2241 : std_logic_vector(63 downto 0);
    signal tmp17_2247 : std_logic_vector(63 downto 0);
    signal tmp18_2253 : std_logic_vector(0 downto 0);
    signal tmp20_1761 : std_logic_vector(31 downto 0);
    signal tmp21_1766 : std_logic_vector(31 downto 0);
    signal tmp22_1770 : std_logic_vector(31 downto 0);
    signal tmp23_1775 : std_logic_vector(31 downto 0);
    signal tmp24_1780 : std_logic_vector(63 downto 0);
    signal tmp25_1786 : std_logic_vector(63 downto 0);
    signal tmp26_1792 : std_logic_vector(0 downto 0);
    signal tmp388_2522 : std_logic_vector(15 downto 0);
    signal tmp389_2622 : std_logic_vector(15 downto 0);
    signal tmp393_2627 : std_logic_vector(15 downto 0);
    signal tmp3_2631 : std_logic_vector(63 downto 0);
    signal tmp406_2199 : std_logic_vector(63 downto 0);
    signal tmp407_2205 : std_logic_vector(0 downto 0);
    signal tmp408_2445 : std_logic_vector(63 downto 0);
    signal tmp415_1735 : std_logic_vector(31 downto 0);
    signal tmp417_1740 : std_logic_vector(31 downto 0);
    signal tmp418_1745 : std_logic_vector(63 downto 0);
    signal tmp419_1751 : std_logic_vector(63 downto 0);
    signal tmp420_1757 : std_logic_vector(0 downto 0);
    signal tmp422_1984 : std_logic_vector(63 downto 0);
    signal tmp4_2637 : std_logic_vector(63 downto 0);
    signal tmp6_2641 : std_logic_vector(63 downto 0);
    signal tmp7_2646 : std_logic_vector(63 downto 0);
    signal tmp9_2209 : std_logic_vector(63 downto 0);
    signal tmp_2057 : std_logic_vector(15 downto 0);
    signal tobool218_2476 : std_logic_vector(0 downto 0);
    signal tobool_2015 : std_logic_vector(0 downto 0);
    signal type_cast_1505_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1530_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1555_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1580_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1605_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1630_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1655_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1680_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1715_wire : std_logic_vector(63 downto 0);
    signal type_cast_1721_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1743_wire : std_logic_vector(63 downto 0);
    signal type_cast_1749_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1778_wire : std_logic_vector(63 downto 0);
    signal type_cast_1784_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1790_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1797_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1806_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1808_wire : std_logic_vector(63 downto 0);
    signal type_cast_1827_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1845_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1863_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1881_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1899_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1917_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1935_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1957_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1976_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1982_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1987_wire : std_logic_vector(63 downto 0);
    signal type_cast_1990_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1999_wire : std_logic_vector(63 downto 0);
    signal type_cast_2002_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2007_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2013_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2026_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2032_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2041_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2043_wire : std_logic_vector(15 downto 0);
    signal type_cast_2048_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2050_wire : std_logic_vector(63 downto 0);
    signal type_cast_2055_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2061_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2079_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2101_wire : std_logic_vector(63 downto 0);
    signal type_cast_2106_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2112_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2118_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2169_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2174_wire : std_logic_vector(63 downto 0);
    signal type_cast_2177_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2184_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2197_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2203_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2239_wire : std_logic_vector(63 downto 0);
    signal type_cast_2245_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2251_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2258_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2267_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2269_wire : std_logic_vector(63 downto 0);
    signal type_cast_2288_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2306_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2324_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2342_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2360_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2378_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2396_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2418_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2437_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2443_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2448_wire : std_logic_vector(63 downto 0);
    signal type_cast_2451_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2460_wire : std_logic_vector(63 downto 0);
    signal type_cast_2463_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2468_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2474_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2487_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2497_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2506_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2508_wire : std_logic_vector(15 downto 0);
    signal type_cast_2513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2515_wire : std_logic_vector(63 downto 0);
    signal type_cast_2520_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2526_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2544_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2566_wire : std_logic_vector(63 downto 0);
    signal type_cast_2571_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2577_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2583_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2620_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2635_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2653_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2655_wire : std_logic_vector(63 downto 0);
    signal type_cast_2671_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2684_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2701_wire : std_logic_vector(63 downto 0);
    signal type_cast_2716_wire : std_logic_vector(63 downto 0);
    signal type_cast_2735_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2750_wire : std_logic_vector(63 downto 0);
    signal type_cast_2753_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2767_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2777_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2787_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2797_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2807_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2817_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2827_wire_constant : std_logic_vector(63 downto 0);
    signal umax19_2260 : std_logic_vector(63 downto 0);
    signal umax27_1799 : std_logic_vector(63 downto 0);
    signal umax421_1978 : std_logic_vector(63 downto 0);
    signal umax_2439 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1814_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1814_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1814_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1814_resized_base_address <= "00000000000000";
    array_obj_ref_2130_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2130_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2130_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2130_resized_base_address <= "00000000000000";
    array_obj_ref_2275_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2275_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2275_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2275_resized_base_address <= "00000000000000";
    array_obj_ref_2595_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2595_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2595_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2595_resized_base_address <= "00000000000000";
    ptr_deref_1951_word_offset_0 <= "00000000000000";
    ptr_deref_2134_word_offset_0 <= "00000000000000";
    ptr_deref_2412_word_offset_0 <= "00000000000000";
    ptr_deref_2599_word_offset_0 <= "00000000000000";
    type_cast_1505_wire_constant <= "00000000000000000000000000001000";
    type_cast_1530_wire_constant <= "0000000000001000";
    type_cast_1555_wire_constant <= "0000000000001000";
    type_cast_1580_wire_constant <= "0000000000001000";
    type_cast_1605_wire_constant <= "0000000000001000";
    type_cast_1630_wire_constant <= "0000000000001000";
    type_cast_1655_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1680_wire_constant <= "0000000000001000";
    type_cast_1721_wire_constant <= "00000000000000000000000000000011";
    type_cast_1749_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1784_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1790_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1797_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1806_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1827_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1845_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1863_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1881_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1899_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1917_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1935_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1957_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1976_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1982_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1990_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2002_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2007_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_2013_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2026_wire_constant <= "00000000000000000000000000000001";
    type_cast_2032_wire_constant <= "00000000000000000000000000000110";
    type_cast_2041_wire_constant <= "0000000000000000";
    type_cast_2048_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2055_wire_constant <= "0000000000000001";
    type_cast_2061_wire_constant <= "0000000000000001";
    type_cast_2079_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2106_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_2112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2118_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2169_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2177_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2184_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_2197_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2203_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2245_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2251_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2258_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2267_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2288_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2306_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2324_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2342_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2360_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2378_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2396_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2418_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2437_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2443_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2451_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2463_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2468_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_2474_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2487_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2497_wire_constant <= "00000000000000000000000000000110";
    type_cast_2506_wire_constant <= "0000000000000000";
    type_cast_2513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2520_wire_constant <= "0000000000000001";
    type_cast_2526_wire_constant <= "0000000000000001";
    type_cast_2544_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2571_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_2577_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2583_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2620_wire_constant <= "1111111111111111";
    type_cast_2635_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2653_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2671_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_2684_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2735_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2753_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2767_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2777_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_2787_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2797_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2807_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2817_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2827_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    phi_stmt_1802: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1806_wire_constant & type_cast_1808_wire;
      req <= phi_stmt_1802_req_0 & phi_stmt_1802_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1802",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1802_ack_0,
          idata => idata,
          odata => indvar425_1802,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1802
    phi_stmt_1996: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1999_wire & type_cast_2002_wire_constant;
      req <= phi_stmt_1996_req_0 & phi_stmt_1996_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1996",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1996_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_1996,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1996
    phi_stmt_2037: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2041_wire_constant & type_cast_2043_wire;
      req <= phi_stmt_2037_req_0 & phi_stmt_2037_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2037",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2037_ack_0,
          idata => idata,
          odata => nx_x022x_xi_2037,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2037
    phi_stmt_2044: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2048_wire_constant & type_cast_2050_wire;
      req <= phi_stmt_2044_req_0 & phi_stmt_2044_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2044",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2044_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_2044,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2044
    phi_stmt_2098: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2101_wire;
      req(0) <= phi_stmt_2098_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2098",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2098_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_2098,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2098
    phi_stmt_2263: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2267_wire_constant & type_cast_2269_wire;
      req <= phi_stmt_2263_req_0 & phi_stmt_2263_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2263",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2263_ack_0,
          idata => idata,
          odata => indvar411_2263,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2263
    phi_stmt_2457: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2460_wire & type_cast_2463_wire_constant;
      req <= phi_stmt_2457_req_0 & phi_stmt_2457_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2457",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2457_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_2457,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2457
    phi_stmt_2502: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2506_wire_constant & type_cast_2508_wire;
      req <= phi_stmt_2502_req_0 & phi_stmt_2502_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2502",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2502_ack_0,
          idata => idata,
          odata => nx_x022x_xi357_2502,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2502
    phi_stmt_2509: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2513_wire_constant & type_cast_2515_wire;
      req <= phi_stmt_2509_req_0 & phi_stmt_2509_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2509",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2509_ack_0,
          idata => idata,
          odata => elementx_x021x_xi358_2509,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2509
    phi_stmt_2563: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2566_wire;
      req(0) <= phi_stmt_2563_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2563",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2563_ack_0,
          idata => idata,
          odata => shl8x_xi362x_xlcssa_2563,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2563
    phi_stmt_2649: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2653_wire_constant & type_cast_2655_wire;
      req <= phi_stmt_2649_req_0 & phi_stmt_2649_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2649",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2649_ack_0,
          idata => idata,
          odata => indvar_2649,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2649
    -- flow-through select operator MUX_1798_inst
    umax27_1799 <= tmp25_1786 when (tmp26_1792(0) /=  '0') else type_cast_1797_wire_constant;
    -- flow-through select operator MUX_1977_inst
    umax421_1978 <= tmp419_1751 when (tmp420_1757(0) /=  '0') else type_cast_1976_wire_constant;
    -- flow-through select operator MUX_2259_inst
    umax19_2260 <= tmp17_2247 when (tmp18_2253(0) /=  '0') else type_cast_2258_wire_constant;
    -- flow-through select operator MUX_2438_inst
    umax_2439 <= tmp406_2199 when (tmp407_2205(0) /=  '0') else type_cast_2437_wire_constant;
    addr_of_1815_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1815_final_reg_req_0;
      addr_of_1815_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1815_final_reg_req_1;
      addr_of_1815_final_reg_ack_1<= rack(0);
      addr_of_1815_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1815_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1814_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1816,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2131_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2131_final_reg_req_0;
      addr_of_2131_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2131_final_reg_req_1;
      addr_of_2131_final_reg_ack_1<= rack(0);
      addr_of_2131_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2131_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2130_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_2132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2276_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2276_final_reg_req_0;
      addr_of_2276_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2276_final_reg_req_1;
      addr_of_2276_final_reg_ack_1<= rack(0);
      addr_of_2276_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2276_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2275_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_2277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2596_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2596_final_reg_req_0;
      addr_of_2596_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2596_final_reg_req_1;
      addr_of_2596_final_reg_ack_1<= rack(0);
      addr_of_2596_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2596_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2595_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_2597,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1500_inst_req_0;
      type_cast_1500_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1500_inst_req_1;
      type_cast_1500_inst_ack_1<= rack(0);
      type_cast_1500_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1500_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_1501,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1513_inst_req_0;
      type_cast_1513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1513_inst_req_1;
      type_cast_1513_inst_ack_1<= rack(0);
      type_cast_1513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1510,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1525_inst_req_0;
      type_cast_1525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1525_inst_req_1;
      type_cast_1525_inst_ack_1<= rack(0);
      type_cast_1525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1522,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_1526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1538_inst_req_0;
      type_cast_1538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1538_inst_req_1;
      type_cast_1538_inst_ack_1<= rack(0);
      type_cast_1538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_1535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1550_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1550_inst_req_0;
      type_cast_1550_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1550_inst_req_1;
      type_cast_1550_inst_ack_1<= rack(0);
      type_cast_1550_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1550_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1547,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_1551,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1563_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1563_inst_req_0;
      type_cast_1563_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1563_inst_req_1;
      type_cast_1563_inst_ack_1<= rack(0);
      type_cast_1563_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1563_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_1560,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1564,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1575_inst_req_0;
      type_cast_1575_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1575_inst_req_1;
      type_cast_1575_inst_ack_1<= rack(0);
      type_cast_1575_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1575_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_1572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1576,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1588_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1588_inst_req_0;
      type_cast_1588_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1588_inst_req_1;
      type_cast_1588_inst_ack_1<= rack(0);
      type_cast_1588_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1588_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_1585,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1589,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1600_inst_req_0;
      type_cast_1600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1600_inst_req_1;
      type_cast_1600_inst_ack_1<= rack(0);
      type_cast_1600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_1597,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1601,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1613_inst_req_0;
      type_cast_1613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1613_inst_req_1;
      type_cast_1613_inst_ack_1<= rack(0);
      type_cast_1613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_1610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_1614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1625_inst_req_0;
      type_cast_1625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1625_inst_req_1;
      type_cast_1625_inst_ack_1<= rack(0);
      type_cast_1625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1625_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_1622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1626,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1638_inst_req_0;
      type_cast_1638_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1638_inst_req_1;
      type_cast_1638_inst_ack_1<= rack(0);
      type_cast_1638_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1638_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_1635,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1639,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1650_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1650_inst_req_0;
      type_cast_1650_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1650_inst_req_1;
      type_cast_1650_inst_ack_1<= rack(0);
      type_cast_1650_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1650_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_1647,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_1651,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1663_inst_req_0;
      type_cast_1663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1663_inst_req_1;
      type_cast_1663_inst_ack_1<= rack(0);
      type_cast_1663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1663_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_1660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1675_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1675_inst_req_0;
      type_cast_1675_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1675_inst_req_1;
      type_cast_1675_inst_ack_1<= rack(0);
      type_cast_1675_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1675_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_1672,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1676,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1688_inst_req_0;
      type_cast_1688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1688_inst_req_1;
      type_cast_1688_inst_ack_1<= rack(0);
      type_cast_1688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_1685,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_1689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1697_inst_req_0;
      type_cast_1697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1697_inst_req_1;
      type_cast_1697_inst_ack_1<= rack(0);
      type_cast_1697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1544,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1701_inst_req_0;
      type_cast_1701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1701_inst_req_1;
      type_cast_1701_inst_ack_1<= rack(0);
      type_cast_1701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1569,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_1702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1716_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1716_inst_req_0;
      type_cast_1716_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1716_inst_req_1;
      type_cast_1716_inst_ack_1<= rack(0);
      type_cast_1716_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1716_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1715_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1717,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1744_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1744_inst_req_0;
      type_cast_1744_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1744_inst_req_1;
      type_cast_1744_inst_ack_1<= rack(0);
      type_cast_1744_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1744_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1743_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp418_1745,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1760_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1760_inst_req_0;
      type_cast_1760_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1760_inst_req_1;
      type_cast_1760_inst_ack_1<= rack(0);
      type_cast_1760_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1760_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1544,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1761,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1769_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1769_inst_req_0;
      type_cast_1769_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1769_inst_req_1;
      type_cast_1769_inst_ack_1<= rack(0);
      type_cast_1769_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1769_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1569,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp22_1770,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1779_inst_req_0;
      type_cast_1779_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1779_inst_req_1;
      type_cast_1779_inst_ack_1<= rack(0);
      type_cast_1779_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1779_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1778_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_1780,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1808_inst_req_0;
      type_cast_1808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1808_inst_req_1;
      type_cast_1808_inst_ack_1<= rack(0);
      type_cast_1808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext426_1959,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1808_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1822_inst_req_0;
      type_cast_1822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1822_inst_req_1;
      type_cast_1822_inst_ack_1<= rack(0);
      type_cast_1822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_1819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1835_inst_req_0;
      type_cast_1835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1835_inst_req_1;
      type_cast_1835_inst_ack_1<= rack(0);
      type_cast_1835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_1832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_1836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1853_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1853_inst_req_0;
      type_cast_1853_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1853_inst_req_1;
      type_cast_1853_inst_ack_1<= rack(0);
      type_cast_1853_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1853_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_1850,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_1854,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1871_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1871_inst_req_0;
      type_cast_1871_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1871_inst_req_1;
      type_cast_1871_inst_ack_1<= rack(0);
      type_cast_1871_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1871_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_1868,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1872,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1889_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1889_inst_req_0;
      type_cast_1889_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1889_inst_req_1;
      type_cast_1889_inst_ack_1<= rack(0);
      type_cast_1889_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1889_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_1886,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_1890,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1907_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1907_inst_req_0;
      type_cast_1907_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1907_inst_req_1;
      type_cast_1907_inst_ack_1<= rack(0);
      type_cast_1907_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1907_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_1904,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_1908,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1925_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1925_inst_req_0;
      type_cast_1925_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1925_inst_req_1;
      type_cast_1925_inst_ack_1<= rack(0);
      type_cast_1925_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1925_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_1922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_1926,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1943_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1943_inst_req_0;
      type_cast_1943_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1943_inst_req_1;
      type_cast_1943_inst_ack_1<= rack(0);
      type_cast_1943_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1943_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_1940,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_1944,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1987_inst
    process(tmp422_1984) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp422_1984(63 downto 0);
      type_cast_1987_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1992_inst
    process(ASHR_i64_i64_1991_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1991_wire(63 downto 0);
      phitmp_1993 <= tmp_var; -- 
    end process;
    type_cast_1999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1999_inst_req_0;
      type_cast_1999_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1999_inst_req_1;
      type_cast_1999_inst_ack_1<= rack(0);
      type_cast_1999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1999_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_1993,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1999_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2043_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2043_inst_req_0;
      type_cast_2043_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2043_inst_req_1;
      type_cast_2043_inst_ack_1<= rack(0);
      type_cast_2043_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2043_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_34_2063,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2043_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2050_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2050_inst_req_0;
      type_cast_2050_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2050_inst_req_1;
      type_cast_2050_inst_ack_1<= rack(0);
      type_cast_2050_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2050_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_2081,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2050_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2069_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2069_inst_req_0;
      type_cast_2069_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2069_inst_req_1;
      type_cast_2069_inst_ack_1<= rack(0);
      type_cast_2069_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2069_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_2066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_2070,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2084_inst_req_0;
      type_cast_2084_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2084_inst_req_1;
      type_cast_2084_inst_ack_1<= rack(0);
      type_cast_2084_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2084_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_2057,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_2085,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2101_inst_req_0;
      type_cast_2101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2101_inst_req_1;
      type_cast_2101_inst_ack_1<= rack(0);
      type_cast_2101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_2081,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2101_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2141_inst_req_0;
      type_cast_2141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2141_inst_req_1;
      type_cast_2141_inst_ack_1<= rack(0);
      type_cast_2141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1569,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_2142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2145_inst_req_0;
      type_cast_2145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2145_inst_req_1;
      type_cast_2145_inst_ack_1<= rack(0);
      type_cast_2145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_1694,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_2146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2149_inst_req_0;
      type_cast_2149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2149_inst_req_1;
      type_cast_2149_inst_ack_1<= rack(0);
      type_cast_2149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_2150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2174_inst
    process(sext_2171) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_2171(63 downto 0);
      type_cast_2174_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2179_inst
    process(ASHR_i64_i64_2178_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_2178_wire(63 downto 0);
      conv155_2180 <= tmp_var; -- 
    end process;
    type_cast_2208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2208_inst_req_0;
      type_cast_2208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2208_inst_req_1;
      type_cast_2208_inst_ack_1<= rack(0);
      type_cast_2208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp9_2209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2217_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2217_inst_req_0;
      type_cast_2217_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2217_inst_req_1;
      type_cast_2217_inst_ack_1<= rack(0);
      type_cast_2217_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2217_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1569,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp11_2218,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2226_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2226_inst_req_0;
      type_cast_2226_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2226_inst_req_1;
      type_cast_2226_inst_ack_1<= rack(0);
      type_cast_2226_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2226_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_1694,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_2227,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2235_inst_req_0;
      type_cast_2235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2235_inst_req_1;
      type_cast_2235_inst_ack_1<= rack(0);
      type_cast_2235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_2232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_2236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2240_inst_req_0;
      type_cast_2240_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2240_inst_req_1;
      type_cast_2240_inst_ack_1<= rack(0);
      type_cast_2240_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2239_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp16_2241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2269_inst_req_0;
      type_cast_2269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2269_inst_req_1;
      type_cast_2269_inst_ack_1<= rack(0);
      type_cast_2269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext412_2420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2269_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2283_inst_req_0;
      type_cast_2283_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2283_inst_req_1;
      type_cast_2283_inst_ack_1<= rack(0);
      type_cast_2283_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2283_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_2280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_2284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2296_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2296_inst_req_0;
      type_cast_2296_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2296_inst_req_1;
      type_cast_2296_inst_ack_1<= rack(0);
      type_cast_2296_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2296_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_2293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_2297,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2314_inst_req_0;
      type_cast_2314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2314_inst_req_1;
      type_cast_2314_inst_ack_1<= rack(0);
      type_cast_2314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_2311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_2315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2332_inst_req_0;
      type_cast_2332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2332_inst_req_1;
      type_cast_2332_inst_ack_1<= rack(0);
      type_cast_2332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_2329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_2333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2350_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2350_inst_req_0;
      type_cast_2350_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2350_inst_req_1;
      type_cast_2350_inst_ack_1<= rack(0);
      type_cast_2350_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2350_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_2347,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_2351,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2368_inst_req_0;
      type_cast_2368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2368_inst_req_1;
      type_cast_2368_inst_ack_1<= rack(0);
      type_cast_2368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_2365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_2369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2386_inst_req_0;
      type_cast_2386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2386_inst_req_1;
      type_cast_2386_inst_ack_1<= rack(0);
      type_cast_2386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_2383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_2387,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2404_inst_req_0;
      type_cast_2404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2404_inst_req_1;
      type_cast_2404_inst_ack_1<= rack(0);
      type_cast_2404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2404_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_2401,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_2405,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2448_inst
    process(tmp408_2445) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp408_2445(63 downto 0);
      type_cast_2448_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2453_inst
    process(ASHR_i64_i64_2452_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_2452_wire(63 downto 0);
      phitmp387_2454 <= tmp_var; -- 
    end process;
    type_cast_2460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2460_inst_req_0;
      type_cast_2460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2460_inst_req_1;
      type_cast_2460_inst_ack_1<= rack(0);
      type_cast_2460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp387_2454,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2460_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2492_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2492_inst_req_0;
      type_cast_2492_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2492_inst_req_1;
      type_cast_2492_inst_ack_1<= rack(0);
      type_cast_2492_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2492_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_56_2489,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi354_2493,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2508_inst_req_0;
      type_cast_2508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2508_inst_req_1;
      type_cast_2508_inst_ack_1<= rack(0);
      type_cast_2508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_68_2528,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2508_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2515_inst_req_0;
      type_cast_2515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2515_inst_req_1;
      type_cast_2515_inst_ack_1<= rack(0);
      type_cast_2515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi362_2546,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2515_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2534_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2534_inst_req_0;
      type_cast_2534_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2534_inst_req_1;
      type_cast_2534_inst_ack_1<= rack(0);
      type_cast_2534_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2534_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi359_2531,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi360_2535,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2549_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2549_inst_req_0;
      type_cast_2549_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2549_inst_req_1;
      type_cast_2549_inst_ack_1<= rack(0);
      type_cast_2549_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2549_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp388_2522,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi363_2550,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2566_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2566_inst_req_0;
      type_cast_2566_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2566_inst_req_1;
      type_cast_2566_inst_ack_1<= rack(0);
      type_cast_2566_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2566_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi362_2546,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2566_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2630_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2630_inst_req_0;
      type_cast_2630_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2630_inst_req_1;
      type_cast_2630_inst_ack_1<= rack(0);
      type_cast_2630_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2630_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp389_2622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_2631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2640_inst_req_0;
      type_cast_2640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2640_inst_req_1;
      type_cast_2640_inst_ack_1<= rack(0);
      type_cast_2640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp393_2627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_2641,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2655_inst_req_0;
      type_cast_2655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2655_inst_req_1;
      type_cast_2655_inst_ack_1<= rack(0);
      type_cast_2655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2686,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2655_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2702_inst_req_0;
      type_cast_2702_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2702_inst_req_1;
      type_cast_2702_inst_ack_1<= rack(0);
      type_cast_2702_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2702_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2701_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_2703,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2717_inst_req_0;
      type_cast_2717_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2717_inst_req_1;
      type_cast_2717_inst_ack_1<= rack(0);
      type_cast_2717_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2717_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2716_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_2718,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2726_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2726_inst_req_0;
      type_cast_2726_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2726_inst_req_1;
      type_cast_2726_inst_ack_1<= rack(0);
      type_cast_2726_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2726_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add43_1619,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv281_2727,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2730_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2730_inst_req_0;
      type_cast_2730_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2730_inst_req_1;
      type_cast_2730_inst_ack_1<= rack(0);
      type_cast_2730_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2730_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_1594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv283_2731,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2750_inst
    process(sext352_2747) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext352_2747(63 downto 0);
      type_cast_2750_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2755_inst
    process(ASHR_i64_i64_2754_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_2754_wire(63 downto 0);
      conv288_2756 <= tmp_var; -- 
    end process;
    type_cast_2762_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2762_inst_req_0;
      type_cast_2762_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2762_inst_req_1;
      type_cast_2762_inst_ack_1<= rack(0);
      type_cast_2762_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2762_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_2723,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv292_2763,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2772_inst_req_0;
      type_cast_2772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2772_inst_req_1;
      type_cast_2772_inst_ack_1<= rack(0);
      type_cast_2772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr295_2769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv298_2773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2782_inst_req_0;
      type_cast_2782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2782_inst_req_1;
      type_cast_2782_inst_ack_1<= rack(0);
      type_cast_2782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr301_2779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_2783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2792_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2792_inst_req_0;
      type_cast_2792_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2792_inst_req_1;
      type_cast_2792_inst_ack_1<= rack(0);
      type_cast_2792_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2792_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr307_2789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv310_2793,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2802_inst_req_0;
      type_cast_2802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2802_inst_req_1;
      type_cast_2802_inst_ack_1<= rack(0);
      type_cast_2802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr313_2799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv316_2803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2812_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2812_inst_req_0;
      type_cast_2812_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2812_inst_req_1;
      type_cast_2812_inst_ack_1<= rack(0);
      type_cast_2812_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2812_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr319_2809,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_2813,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2822_inst_req_0;
      type_cast_2822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2822_inst_req_1;
      type_cast_2822_inst_ack_1<= rack(0);
      type_cast_2822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr325_2819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv328_2823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2832_inst_req_0;
      type_cast_2832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2832_inst_req_1;
      type_cast_2832_inst_ack_1<= rack(0);
      type_cast_2832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr331_2829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv334_2833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1814_index_1_rename
    process(R_indvar425_1813_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar425_1813_resized;
      ov(13 downto 0) := iv;
      R_indvar425_1813_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1814_index_1_resize
    process(indvar425_1802) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar425_1802;
      ov := iv(13 downto 0);
      R_indvar425_1813_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1814_root_address_inst
    process(array_obj_ref_1814_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1814_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1814_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2130_index_1_rename
    process(R_ix_x0x_xlcssa_2129_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_2129_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_2129_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2130_index_1_resize
    process(ix_x0x_xlcssa_1996) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_1996;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_2129_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2130_root_address_inst
    process(array_obj_ref_2130_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2130_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2130_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2275_index_1_rename
    process(R_indvar411_2274_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar411_2274_resized;
      ov(13 downto 0) := iv;
      R_indvar411_2274_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2275_index_1_resize
    process(indvar411_2263) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar411_2263;
      ov := iv(13 downto 0);
      R_indvar411_2274_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2275_root_address_inst
    process(array_obj_ref_2275_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2275_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2275_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2595_index_1_rename
    process(R_ix_x1x_xlcssa_2594_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_2594_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_2594_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2595_index_1_resize
    process(ix_x1x_xlcssa_2457) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_2457;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_2594_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2595_root_address_inst
    process(array_obj_ref_2595_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2595_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2595_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1951_addr_0
    process(ptr_deref_1951_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1951_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1951_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1951_base_resize
    process(arrayidx_1816) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1816;
      ov := iv(13 downto 0);
      ptr_deref_1951_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1951_gather_scatter
    process(add132_1949) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_1949;
      ov(63 downto 0) := iv;
      ptr_deref_1951_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1951_root_address_inst
    process(ptr_deref_1951_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1951_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1951_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2134_addr_0
    process(ptr_deref_2134_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2134_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2134_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2134_base_resize
    process(arrayidx143_2132) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_2132;
      ov := iv(13 downto 0);
      ptr_deref_2134_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2134_gather_scatter
    process(shl14x_xi_2125) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_2125;
      ov(63 downto 0) := iv;
      ptr_deref_2134_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2134_root_address_inst
    process(ptr_deref_2134_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2134_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2134_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2412_addr_0
    process(ptr_deref_2412_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2412_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2412_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2412_base_resize
    process(arrayidx211_2277) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_2277;
      ov := iv(13 downto 0);
      ptr_deref_2412_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2412_gather_scatter
    process(add207_2410) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_2410;
      ov(63 downto 0) := iv;
      ptr_deref_2412_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2412_root_address_inst
    process(ptr_deref_2412_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2412_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2412_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2599_addr_0
    process(ptr_deref_2599_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2599_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2599_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2599_base_resize
    process(arrayidx226_2597) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_2597;
      ov := iv(13 downto 0);
      ptr_deref_2599_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2599_gather_scatter
    process(shl14x_xi372_2590) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi372_2590;
      ov(63 downto 0) := iv;
      ptr_deref_2599_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2599_root_address_inst
    process(ptr_deref_2599_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2599_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2599_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1724_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp383_1723;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1724_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1724_branch_req_0,
          ack0 => if_stmt_1724_branch_ack_0,
          ack1 => if_stmt_1724_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1965_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond28_1964;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1965_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1965_branch_req_0,
          ack0 => if_stmt_1965_branch_ack_0,
          ack1 => if_stmt_1965_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2016_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_2015;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2016_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2016_branch_req_0,
          ack0 => if_stmt_2016_branch_ack_0,
          ack1 => if_stmt_2016_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2091_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_2090;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2091_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2091_branch_req_0,
          ack0 => if_stmt_2091_branch_ack_0,
          ack1 => if_stmt_2091_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2187_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161379_2186;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2187_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2187_branch_req_0,
          ack0 => if_stmt_2187_branch_ack_0,
          ack1 => if_stmt_2187_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2426_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_2425;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2426_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2426_branch_req_0,
          ack0 => if_stmt_2426_branch_ack_0,
          ack1 => if_stmt_2426_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2477_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_2476;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2477_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2477_branch_req_0,
          ack0 => if_stmt_2477_branch_ack_0,
          ack1 => if_stmt_2477_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2556_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi364_2555;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2556_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2556_branch_req_0,
          ack0 => if_stmt_2556_branch_ack_0,
          ack1 => if_stmt_2556_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2692_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_2691;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2692_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2692_branch_req_0,
          ack0 => if_stmt_2692_branch_ack_0,
          ack1 => if_stmt_2692_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2056_inst
    process(nx_x022x_xi_2037) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_2037, type_cast_2055_wire_constant, tmp_var);
      tmp_2057 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2062_inst
    process(nx_x022x_xi_2037) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_2037, type_cast_2061_wire_constant, tmp_var);
      iNsTr_34_2063 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2521_inst
    process(nx_x022x_xi357_2502) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi357_2502, type_cast_2520_wire_constant, tmp_var);
      tmp388_2522 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2527_inst
    process(nx_x022x_xi357_2502) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi357_2502, type_cast_2526_wire_constant, tmp_var);
      iNsTr_68_2528 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2621_inst
    process(add53_1644) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_1644, type_cast_2620_wire_constant, tmp_var);
      tmp389_2622 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1958_inst
    process(indvar425_1802) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar425_1802, type_cast_1957_wire_constant, tmp_var);
      indvarx_xnext426_1959 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2419_inst
    process(indvar411_2263) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar411_2263, type_cast_2418_wire_constant, tmp_var);
      indvarx_xnext412_2420 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2636_inst
    process(tmp3_2631) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2631, type_cast_2635_wire_constant, tmp_var);
      tmp4_2637 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2685_inst
    process(indvar_2649) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2649, type_cast_2684_wire_constant, tmp_var);
      indvarx_xnext_2686 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2033_inst
    process(conv2x_xi_2028) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_2028, type_cast_2032_wire_constant, tmp_var);
      shlx_xi_2034 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2498_inst
    process(conv2x_xi354_2493) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi354_2493, type_cast_2497_wire_constant, tmp_var);
      shlx_xi355_2499 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2008_inst
    process(conv83_1717) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_1717, type_cast_2007_wire_constant, tmp_var);
      and_2009 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2113_inst
    process(Bx_xnot_2108) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_2108, type_cast_2112_wire_constant, tmp_var);
      add1216x_xi_2114 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2469_inst
    process(conv155_2180) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_2180, type_cast_2468_wire_constant, tmp_var);
      and217_2470 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2578_inst
    process(iNsTr_94_2573) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_94_2573, type_cast_2577_wire_constant, tmp_var);
      add1216x_xi370_2579 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2672_inst
    process(mul253_2661) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul253_2661, type_cast_2671_wire_constant, tmp_var);
      conv254_2673 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1991_inst
    process(type_cast_1987_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1987_wire, type_cast_1990_wire_constant, tmp_var);
      ASHR_i64_i64_1991_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_2178_inst
    process(type_cast_2174_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2174_wire, type_cast_2177_wire_constant, tmp_var);
      ASHR_i64_i64_2178_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_2452_inst
    process(type_cast_2448_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2448_wire, type_cast_2451_wire_constant, tmp_var);
      ASHR_i64_i64_2452_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_2754_inst
    process(type_cast_2750_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2750_wire, type_cast_2753_wire_constant, tmp_var);
      ASHR_i64_i64_2754_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1963_inst
    process(indvarx_xnext426_1959, umax27_1799) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext426_1959, umax27_1799, tmp_var);
      exitcond28_1964 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2014_inst
    process(and_2009) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_2009, type_cast_2013_wire_constant, tmp_var);
      tobool_2015 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2424_inst
    process(indvarx_xnext412_2420, umax19_2260) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext412_2420, umax19_2260, tmp_var);
      exitcond_2425 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2475_inst
    process(and217_2470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_2470, type_cast_2474_wire_constant, tmp_var);
      tobool218_2476 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2690_inst
    process(indvarx_xnext_2686, tmp4_2637) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_2686, tmp4_2637, tmp_var);
      exitcond5_2691 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1750_inst
    process(tmp418_1745) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp418_1745, type_cast_1749_wire_constant, tmp_var);
      tmp419_1751 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1785_inst
    process(tmp24_1780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp24_1780, type_cast_1784_wire_constant, tmp_var);
      tmp25_1786 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2198_inst
    process(conv155_2180) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_2180, type_cast_2197_wire_constant, tmp_var);
      tmp406_2199 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2246_inst
    process(tmp16_2241) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp16_2241, type_cast_2245_wire_constant, tmp_var);
      tmp17_2247 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2768_inst
    process(sub_2723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2723, type_cast_2767_wire_constant, tmp_var);
      shr295_2769 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2778_inst
    process(sub_2723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2723, type_cast_2777_wire_constant, tmp_var);
      shr301_2779 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2788_inst
    process(sub_2723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2723, type_cast_2787_wire_constant, tmp_var);
      shr307_2789 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2798_inst
    process(sub_2723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2723, type_cast_2797_wire_constant, tmp_var);
      shr313_2799 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2808_inst
    process(sub_2723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2723, type_cast_2807_wire_constant, tmp_var);
      shr319_2809 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2818_inst
    process(sub_2723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2723, type_cast_2817_wire_constant, tmp_var);
      shr325_2819 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2828_inst
    process(sub_2723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2723, type_cast_2827_wire_constant, tmp_var);
      shr331_2829 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2626_inst
    process(add73_1694, add23_1569) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1694, add23_1569, tmp_var);
      tmp393_2627 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1706_inst
    process(conv79_1698, add_1519) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_1698, add_1519, tmp_var);
      mul_1707 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1711_inst
    process(mul_1707, conv81_1702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1707, conv81_1702, tmp_var);
      mul82_1712 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1734_inst
    process(add_1519, conv79_1698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1519, conv79_1698, tmp_var);
      tmp415_1735 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1739_inst
    process(tmp415_1735, conv81_1702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp415_1735, conv81_1702, tmp_var);
      tmp417_1740 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1765_inst
    process(add_1519, tmp20_1761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1519, tmp20_1761, tmp_var);
      tmp21_1766 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1774_inst
    process(tmp21_1766, tmp22_1770) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp21_1766, tmp22_1770, tmp_var);
      tmp23_1775 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2154_inst
    process(conv153_2150, conv145_2142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_2150, conv145_2142, tmp_var);
      mul148_2155 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2159_inst
    process(mul148_2155, add63_1669) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_2155, add63_1669, tmp_var);
      mul151_2160 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2164_inst
    process(mul151_2160, conv147_2146) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_2160, conv147_2146, tmp_var);
      mul154_2165 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2213_inst
    process(add63_1669, tmp9_2209) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_1669, tmp9_2209, tmp_var);
      tmp10_2214 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2222_inst
    process(tmp10_2214, tmp11_2218) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp10_2214, tmp11_2218, tmp_var);
      tmp12_2223 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2231_inst
    process(tmp12_2223, tmp13_2227) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_2223, tmp13_2227, tmp_var);
      tmp14_2232 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2645_inst
    process(add63_1669, tmp6_2641) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_1669, tmp6_2641, tmp_var);
      tmp7_2646 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2660_inst
    process(tmp7_2646, indvar_2649) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp7_2646, indvar_2649, tmp_var);
      mul253_2661 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2741_inst
    process(mul284_2737, conv281_2727) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul284_2737, conv281_2727, tmp_var);
      mul287_2742 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2746_inst
    process(mul287_2742, conv153_2150) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul287_2742, conv153_2150, tmp_var);
      sext352_2747 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1543_inst
    process(shl10_1532, conv12_1539) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_1532, conv12_1539, tmp_var);
      add13_1544 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1568_inst
    process(shl20_1557, conv22_1564) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_1557, conv22_1564, tmp_var);
      add23_1569 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1593_inst
    process(shl30_1582, conv32_1589) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_1582, conv32_1589, tmp_var);
      add33_1594 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1618_inst
    process(shl40_1607, conv42_1614) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_1607, conv42_1614, tmp_var);
      add43_1619 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1643_inst
    process(shl50_1632, conv52_1639) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_1632, conv52_1639, tmp_var);
      add53_1644 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1693_inst
    process(shl70_1682, conv72_1689) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_1682, conv72_1689, tmp_var);
      add73_1694 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1518_inst
    process(shl_1507, conv3_1514) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1507, conv3_1514, tmp_var);
      add_1519 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1668_inst
    process(shl60_1657, conv62_1664) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_1657, conv62_1664, tmp_var);
      add63_1669 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1840_inst
    process(shl92_1829, conv95_1836) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_1829, conv95_1836, tmp_var);
      add96_1841 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1858_inst
    process(shl98_1847, conv101_1854) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_1847, conv101_1854, tmp_var);
      add102_1859 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1876_inst
    process(shl104_1865, conv107_1872) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_1865, conv107_1872, tmp_var);
      add108_1877 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1894_inst
    process(shl110_1883, conv113_1890) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_1883, conv113_1890, tmp_var);
      add114_1895 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1912_inst
    process(shl116_1901, conv119_1908) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_1901, conv119_1908, tmp_var);
      add120_1913 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1930_inst
    process(shl122_1919, conv125_1926) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_1919, conv125_1926, tmp_var);
      add126_1931 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1948_inst
    process(shl128_1937, conv131_1944) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_1937, conv131_1944, tmp_var);
      add132_1949 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2074_inst
    process(conv5x_xi_2070, elementx_x021x_xi_2044) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_2070, elementx_x021x_xi_2044, tmp_var);
      addx_xi_2075 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2301_inst
    process(shl167_2290, conv170_2297) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_2290, conv170_2297, tmp_var);
      add171_2302 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2319_inst
    process(shl173_2308, conv176_2315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_2308, conv176_2315, tmp_var);
      add177_2320 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2337_inst
    process(shl179_2326, conv182_2333) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_2326, conv182_2333, tmp_var);
      add183_2338 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2355_inst
    process(shl185_2344, conv188_2351) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_2344, conv188_2351, tmp_var);
      add189_2356 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2373_inst
    process(shl191_2362, conv194_2369) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_2362, conv194_2369, tmp_var);
      add195_2374 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2391_inst
    process(shl197_2380, conv200_2387) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_2380, conv200_2387, tmp_var);
      add201_2392 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2409_inst
    process(shl203_2398, conv206_2405) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_2398, conv206_2405, tmp_var);
      add207_2410 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2539_inst
    process(conv5x_xi360_2535, elementx_x021x_xi358_2509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi360_2535, elementx_x021x_xi358_2509, tmp_var);
      addx_xi361_2540 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1531_inst
    process(conv9_1526) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_1526, type_cast_1530_wire_constant, tmp_var);
      shl10_1532 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1556_inst
    process(conv19_1551) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_1551, type_cast_1555_wire_constant, tmp_var);
      shl20_1557 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1581_inst
    process(conv29_1576) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_1576, type_cast_1580_wire_constant, tmp_var);
      shl30_1582 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1606_inst
    process(conv39_1601) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_1601, type_cast_1605_wire_constant, tmp_var);
      shl40_1607 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1631_inst
    process(conv49_1626) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1626, type_cast_1630_wire_constant, tmp_var);
      shl50_1632 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1681_inst
    process(conv69_1676) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_1676, type_cast_1680_wire_constant, tmp_var);
      shl70_1682 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1506_inst
    process(conv1_1501) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_1501, type_cast_1505_wire_constant, tmp_var);
      shl_1507 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2027_inst
    process(mul82_1712) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_1712, type_cast_2026_wire_constant, tmp_var);
      conv2x_xi_2028 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1656_inst
    process(conv59_1651) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_1651, type_cast_1655_wire_constant, tmp_var);
      shl60_1657 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1828_inst
    process(conv90_1823) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_1823, type_cast_1827_wire_constant, tmp_var);
      shl92_1829 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1846_inst
    process(add96_1841) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_1841, type_cast_1845_wire_constant, tmp_var);
      shl98_1847 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1864_inst
    process(add102_1859) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_1859, type_cast_1863_wire_constant, tmp_var);
      shl104_1865 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1882_inst
    process(add108_1877) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_1877, type_cast_1881_wire_constant, tmp_var);
      shl110_1883 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1900_inst
    process(add114_1895) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_1895, type_cast_1899_wire_constant, tmp_var);
      shl116_1901 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1918_inst
    process(add120_1913) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_1913, type_cast_1917_wire_constant, tmp_var);
      shl122_1919 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1936_inst
    process(add126_1931) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_1931, type_cast_1935_wire_constant, tmp_var);
      shl128_1937 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1983_inst
    process(umax421_1978) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax421_1978, type_cast_1982_wire_constant, tmp_var);
      tmp422_1984 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2080_inst
    process(addx_xi_2075) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_2075, type_cast_2079_wire_constant, tmp_var);
      shl8x_xi_2081 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2107_inst
    process(conv83_1717) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_1717, type_cast_2106_wire_constant, tmp_var);
      Bx_xnot_2108 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2124_inst
    process(shl8x_xix_xlcssa_2098, sh_promx_xi_2120) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_2098, sh_promx_xi_2120, tmp_var);
      shl14x_xi_2125 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2170_inst
    process(mul154_2165) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_2165, type_cast_2169_wire_constant, tmp_var);
      sext_2171 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2289_inst
    process(conv165_2284) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_2284, type_cast_2288_wire_constant, tmp_var);
      shl167_2290 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2307_inst
    process(add171_2302) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_2302, type_cast_2306_wire_constant, tmp_var);
      shl173_2308 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2325_inst
    process(add177_2320) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_2320, type_cast_2324_wire_constant, tmp_var);
      shl179_2326 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2343_inst
    process(add183_2338) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_2338, type_cast_2342_wire_constant, tmp_var);
      shl185_2344 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2361_inst
    process(add189_2356) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_2356, type_cast_2360_wire_constant, tmp_var);
      shl191_2362 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2379_inst
    process(add195_2374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_2374, type_cast_2378_wire_constant, tmp_var);
      shl197_2380 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2397_inst
    process(add201_2392) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_2392, type_cast_2396_wire_constant, tmp_var);
      shl203_2398 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2444_inst
    process(umax_2439) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_2439, type_cast_2443_wire_constant, tmp_var);
      tmp408_2445 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2488_inst
    process(mul154_2165) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_2165, type_cast_2487_wire_constant, tmp_var);
      iNsTr_56_2489 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2545_inst
    process(addx_xi361_2540) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi361_2540, type_cast_2544_wire_constant, tmp_var);
      shl8x_xi362_2546 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2572_inst
    process(mul154_2165) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_2165, type_cast_2571_wire_constant, tmp_var);
      iNsTr_94_2573 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2589_inst
    process(shl8x_xi362x_xlcssa_2563, sh_promx_xi371_2585) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi362x_xlcssa_2563, sh_promx_xi371_2585, tmp_var);
      shl14x_xi372_2590 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2736_inst
    process(conv283_2731) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv283_2731, type_cast_2735_wire_constant, tmp_var);
      mul284_2737 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_2722_inst
    process(conv276_2718, conv230_2703) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv276_2718, conv230_2703, tmp_var);
      sub_2723 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1722_inst
    process(mul82_1712) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_1712, type_cast_1721_wire_constant, tmp_var);
      cmp383_1723 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1756_inst
    process(tmp419_1751) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp419_1751, type_cast_1755_wire_constant, tmp_var);
      tmp420_1757 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1791_inst
    process(tmp25_1786) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp25_1786, type_cast_1790_wire_constant, tmp_var);
      tmp26_1792 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_2185_inst
    process(conv155_2180) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_2180, type_cast_2184_wire_constant, tmp_var);
      cmp161379_2186 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_2204_inst
    process(tmp406_2199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp406_2199, type_cast_2203_wire_constant, tmp_var);
      tmp407_2205 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_2252_inst
    process(tmp17_2247) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp17_2247, type_cast_2251_wire_constant, tmp_var);
      tmp18_2253 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2089_inst
    process(convx_xi_2085, shlx_xi_2034) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_2085, shlx_xi_2034, tmp_var);
      cmpx_xi_2090 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2554_inst
    process(convx_xi363_2550, shlx_xi355_2499) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi363_2550, shlx_xi355_2499, tmp_var);
      cmpx_xi364_2555 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_2119_inst
    process(add1216x_xi_2114) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_2114, type_cast_2118_wire_constant, tmp_var);
      sh_promx_xi_2120 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_2584_inst
    process(add1216x_xi370_2579) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi370_2579, type_cast_2583_wire_constant, tmp_var);
      sh_promx_xi371_2585 <= tmp_var; --
    end process;
    -- shared split operator group (122) : array_obj_ref_1814_index_offset 
    ApIntAdd_group_122: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar425_1813_scaled;
      array_obj_ref_1814_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1814_index_offset_req_0;
      array_obj_ref_1814_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1814_index_offset_req_1;
      array_obj_ref_1814_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_122_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_122_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- shared split operator group (123) : array_obj_ref_2130_index_offset 
    ApIntAdd_group_123: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_2129_scaled;
      array_obj_ref_2130_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2130_index_offset_req_0;
      array_obj_ref_2130_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2130_index_offset_req_1;
      array_obj_ref_2130_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_123_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_123_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : array_obj_ref_2275_index_offset 
    ApIntAdd_group_124: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar411_2274_scaled;
      array_obj_ref_2275_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2275_index_offset_req_0;
      array_obj_ref_2275_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2275_index_offset_req_1;
      array_obj_ref_2275_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_124_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_124_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : array_obj_ref_2595_index_offset 
    ApIntAdd_group_125: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_2594_scaled;
      array_obj_ref_2595_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2595_index_offset_req_0;
      array_obj_ref_2595_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2595_index_offset_req_1;
      array_obj_ref_2595_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_125_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_125_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- unary operator type_cast_1715_inst
    process(mul82_1712) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_1712, tmp_var);
      type_cast_1715_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1743_inst
    process(tmp417_1740) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp417_1740, tmp_var);
      type_cast_1743_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1778_inst
    process(tmp23_1775) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp23_1775, tmp_var);
      type_cast_1778_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2239_inst
    process(tmp15_2236) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp15_2236, tmp_var);
      type_cast_2239_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2701_inst
    process(call229_2606) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_2606, tmp_var);
      type_cast_2701_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2716_inst
    process(call275_2713) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_2713, tmp_var);
      type_cast_2716_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1951_store_0 ptr_deref_2134_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1951_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2134_store_0_req_0;
      ptr_deref_1951_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2134_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1951_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2134_store_0_req_1;
      ptr_deref_1951_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2134_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1951_word_address_0 & ptr_deref_2134_word_address_0;
      data_in <= ptr_deref_1951_data_0 & ptr_deref_2134_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_2412_store_0 ptr_deref_2599_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2412_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2599_store_0_req_0;
      ptr_deref_2412_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2599_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2412_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2599_store_0_req_1;
      ptr_deref_2412_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2599_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2412_word_address_0 & ptr_deref_2599_word_address_0;
      data_in <= ptr_deref_2412_data_0 & ptr_deref_2599_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_input_done_pipe_2705_inst RPIPE_input_done_pipe_2709_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_input_done_pipe_2705_inst_req_0;
      reqL_unguarded(0) <= RPIPE_input_done_pipe_2709_inst_req_0;
      RPIPE_input_done_pipe_2705_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_input_done_pipe_2709_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_input_done_pipe_2705_inst_req_1;
      reqR_unguarded(0) <= RPIPE_input_done_pipe_2709_inst_req_1;
      RPIPE_input_done_pipe_2705_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_input_done_pipe_2709_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      call270_2706 <= data_out(15 downto 8);
      call273_2710 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_maxpool_input_pipe_1496_inst RPIPE_maxpool_input_pipe_1509_inst RPIPE_maxpool_input_pipe_1521_inst RPIPE_maxpool_input_pipe_1534_inst RPIPE_maxpool_input_pipe_1546_inst RPIPE_maxpool_input_pipe_1559_inst RPIPE_maxpool_input_pipe_1571_inst RPIPE_maxpool_input_pipe_1584_inst RPIPE_maxpool_input_pipe_1596_inst RPIPE_maxpool_input_pipe_1609_inst RPIPE_maxpool_input_pipe_1621_inst RPIPE_maxpool_input_pipe_1634_inst RPIPE_maxpool_input_pipe_1646_inst RPIPE_maxpool_input_pipe_1659_inst RPIPE_maxpool_input_pipe_1671_inst RPIPE_maxpool_input_pipe_1684_inst RPIPE_maxpool_input_pipe_1818_inst RPIPE_maxpool_input_pipe_1831_inst RPIPE_maxpool_input_pipe_1849_inst RPIPE_maxpool_input_pipe_1867_inst RPIPE_maxpool_input_pipe_1885_inst RPIPE_maxpool_input_pipe_1903_inst RPIPE_maxpool_input_pipe_1921_inst RPIPE_maxpool_input_pipe_1939_inst RPIPE_maxpool_input_pipe_2065_inst RPIPE_maxpool_input_pipe_2279_inst RPIPE_maxpool_input_pipe_2292_inst RPIPE_maxpool_input_pipe_2310_inst RPIPE_maxpool_input_pipe_2328_inst RPIPE_maxpool_input_pipe_2346_inst RPIPE_maxpool_input_pipe_2364_inst RPIPE_maxpool_input_pipe_2382_inst RPIPE_maxpool_input_pipe_2400_inst RPIPE_maxpool_input_pipe_2530_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_1496_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_1509_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_1521_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_1534_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_1546_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_1559_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_1571_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_1584_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_1596_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_1609_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_1621_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_1634_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_1646_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_1659_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_1671_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_1684_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_1818_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_1831_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_1849_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_1867_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_1885_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_1903_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1921_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1939_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_2065_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_2279_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_2292_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_2310_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_2328_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_2346_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_2364_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_2382_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_2400_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_2530_inst_req_0;
      RPIPE_maxpool_input_pipe_1496_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_1509_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_1521_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_1534_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_1546_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_1559_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_1571_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_1584_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_1596_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_1609_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_1621_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_1634_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_1646_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_1659_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_1671_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_1684_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_1818_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_1831_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_1849_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_1867_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_1885_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_1903_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_1921_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1939_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_2065_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_2279_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_2292_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_2310_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_2328_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_2346_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_2364_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_2382_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_2400_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_2530_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_1496_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_1509_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_1521_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_1534_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_1546_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_1559_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_1571_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_1584_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_1596_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_1609_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_1621_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_1634_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_1646_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_1659_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_1671_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_1684_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_1818_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_1831_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_1849_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_1867_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_1885_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_1903_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1921_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1939_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_2065_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_2279_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_2292_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_2310_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_2328_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_2346_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_2364_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_2382_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_2400_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_2530_inst_req_1;
      RPIPE_maxpool_input_pipe_1496_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_1509_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_1521_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_1534_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_1546_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_1559_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_1571_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_1584_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_1596_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_1609_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_1621_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_1634_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_1646_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_1659_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_1671_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_1684_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_1818_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_1831_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_1849_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_1867_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_1885_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_1903_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_1921_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1939_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_2065_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_2279_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_2292_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_2310_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_2328_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_2346_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_2364_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_2382_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_2400_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_2530_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call_1497 <= data_out(271 downto 264);
      call2_1510 <= data_out(263 downto 256);
      call6_1522 <= data_out(255 downto 248);
      call11_1535 <= data_out(247 downto 240);
      call16_1547 <= data_out(239 downto 232);
      call21_1560 <= data_out(231 downto 224);
      call26_1572 <= data_out(223 downto 216);
      call31_1585 <= data_out(215 downto 208);
      call36_1597 <= data_out(207 downto 200);
      call41_1610 <= data_out(199 downto 192);
      call46_1622 <= data_out(191 downto 184);
      call51_1635 <= data_out(183 downto 176);
      call56_1647 <= data_out(175 downto 168);
      call61_1660 <= data_out(167 downto 160);
      call66_1672 <= data_out(159 downto 152);
      call71_1685 <= data_out(151 downto 144);
      call89_1819 <= data_out(143 downto 136);
      call93_1832 <= data_out(135 downto 128);
      call99_1850 <= data_out(127 downto 120);
      call105_1868 <= data_out(119 downto 112);
      call111_1886 <= data_out(111 downto 104);
      call117_1904 <= data_out(103 downto 96);
      call123_1922 <= data_out(95 downto 88);
      call129_1940 <= data_out(87 downto 80);
      callx_xi_2066 <= data_out(79 downto 72);
      call164_2280 <= data_out(71 downto 64);
      call168_2293 <= data_out(63 downto 56);
      call174_2311 <= data_out(55 downto 48);
      call180_2329 <= data_out(47 downto 40);
      call186_2347 <= data_out(39 downto 32);
      call192_2365 <= data_out(31 downto 24);
      call198_2383 <= data_out(23 downto 16);
      call204_2401 <= data_out(15 downto 8);
      callx_xi359_2531 <= data_out(7 downto 0);
      maxpool_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_1_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_1", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_2834_inst WPIPE_maxpool_output_pipe_2837_inst WPIPE_maxpool_output_pipe_2840_inst WPIPE_maxpool_output_pipe_2843_inst WPIPE_maxpool_output_pipe_2846_inst WPIPE_maxpool_output_pipe_2849_inst WPIPE_maxpool_output_pipe_2852_inst WPIPE_maxpool_output_pipe_2855_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_2834_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_2837_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_2840_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_2843_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_2846_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_2849_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2852_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2855_inst_req_0;
      WPIPE_maxpool_output_pipe_2834_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_2837_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_2840_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_2843_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_2846_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_2849_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_2852_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2855_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_2834_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_2837_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_2840_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_2843_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_2846_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_2849_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2852_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2855_inst_req_1;
      WPIPE_maxpool_output_pipe_2834_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_2837_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_2840_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_2843_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_2846_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_2849_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_2852_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2855_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv334_2833 & conv328_2823 & conv322_2813 & conv316_2803 & conv310_2793 & conv304_2783 & conv298_2773 & conv292_2763;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_num_out_pipe_2662_inst WPIPE_num_out_pipe_2665_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_num_out_pipe_2662_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_2665_inst_req_0;
      WPIPE_num_out_pipe_2662_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_num_out_pipe_2665_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_num_out_pipe_2662_inst_req_1;
      update_req_unguarded(0) <= WPIPE_num_out_pipe_2665_inst_req_1;
      WPIPE_num_out_pipe_2662_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_num_out_pipe_2665_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= add33_1594 & add43_1619;
      num_out_pipe_write_1_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_output_pipe_2607_inst WPIPE_output_pipe_2610_inst WPIPE_output_pipe_2613_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal sample_req, sample_ack : BooleanArray( 2 downto 0);
      signal update_req, update_ack : BooleanArray( 2 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 2 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      sample_req_unguarded(2) <= WPIPE_output_pipe_2607_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_output_pipe_2610_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_output_pipe_2613_inst_req_0;
      WPIPE_output_pipe_2607_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_output_pipe_2610_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_output_pipe_2613_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(2) <= WPIPE_output_pipe_2607_inst_req_1;
      update_req_unguarded(1) <= WPIPE_output_pipe_2610_inst_req_1;
      update_req_unguarded(0) <= WPIPE_output_pipe_2613_inst_req_1;
      WPIPE_output_pipe_2607_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_output_pipe_2610_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_output_pipe_2613_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      data_in <= add33_1594 & add43_1619 & add53_1644;
      output_pipe_write_2_gI: SplitGuardInterface generic map(name => "output_pipe_write_2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 3, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_2606_call call_stmt_2713_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_2606_call_req_0;
      reqL_unguarded(0) <= call_stmt_2713_call_req_0;
      call_stmt_2606_call_ack_0 <= ackL_unguarded(1);
      call_stmt_2713_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_2606_call_req_1;
      reqR_unguarded(0) <= call_stmt_2713_call_req_1;
      call_stmt_2606_call_ack_1 <= ackR_unguarded(1);
      call_stmt_2713_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call229_2606 <= data_out(127 downto 64);
      call275_2713 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2676_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2676_call_req_0;
      call_stmt_2676_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2676_call_req_1;
      call_stmt_2676_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv254_2673 & add23_1569;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(79 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2680_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2680_call_req_0;
      call_stmt_2680_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2680_call_req_1;
      call_stmt_2680_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add33_1594 & add23_1569 & add13_1544;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 48,
        owidth => 48,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(47 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_2758_call 
    sendB_call_group_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2758_call_req_0;
      call_stmt_2758_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2758_call_req_1;
      call_stmt_2758_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_3_gI: SplitGuardInterface generic map(name => "sendB_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv288_2756;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(63 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe4_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe4_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_6745_start: Boolean;
  signal convolve_CP_6745_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_size_pipe_2883_inst_req_0 : boolean;
  signal RPIPE_size_pipe_2883_inst_req_1 : boolean;
  signal nacc1_3293_2894_buf_req_1 : boolean;
  signal W_store_kernel_3131_delayed_1_0_3233_inst_req_1 : boolean;
  signal SUB_u16_u16_2880_inst_ack_1 : boolean;
  signal W_read_k_3004_delayed_1_0_3084_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_2873_inst_req_1 : boolean;
  signal W_store_kernel_3127_delayed_1_0_3226_inst_ack_1 : boolean;
  signal RPIPE_num_out_pipe_2873_inst_ack_0 : boolean;
  signal W_read_k_3010_delayed_1_0_3093_inst_req_1 : boolean;
  signal phi_stmt_2889_req_0 : boolean;
  signal nacc2_3302_2899_buf_req_0 : boolean;
  signal RPIPE_size_pipe_2883_inst_ack_0 : boolean;
  signal SUB_u16_u16_2880_inst_req_1 : boolean;
  signal SUB_u16_u16_2880_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2873_inst_req_0 : boolean;
  signal SUB_u16_u16_2880_inst_req_0 : boolean;
  signal phi_stmt_2889_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2873_inst_ack_1 : boolean;
  signal W_read_k_3004_delayed_1_0_3084_inst_req_1 : boolean;
  signal phi_stmt_2889_req_1 : boolean;
  signal SUB_u16_u16_2875_inst_ack_1 : boolean;
  signal SUB_u16_u16_2875_inst_req_1 : boolean;
  signal W_store_kernel_3127_delayed_1_0_3226_inst_req_0 : boolean;
  signal W_read_k_3010_delayed_1_0_3093_inst_req_0 : boolean;
  signal SUB_u16_u16_2885_inst_ack_1 : boolean;
  signal SUB_u16_u16_3208_inst_req_0 : boolean;
  signal phi_stmt_2895_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2878_inst_ack_1 : boolean;
  signal W_read_k_3004_delayed_1_0_3084_inst_ack_1 : boolean;
  signal SUB_u16_u16_2885_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_2878_inst_req_1 : boolean;
  signal SUB_u16_u16_3208_inst_req_1 : boolean;
  signal SUB_u16_u16_3208_inst_ack_1 : boolean;
  signal W_read_k_3010_delayed_1_0_3093_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2878_inst_ack_0 : boolean;
  signal nacc1_3293_2894_buf_ack_1 : boolean;
  signal RPIPE_num_out_pipe_2878_inst_req_0 : boolean;
  signal n_col_3276_2909_buf_req_0 : boolean;
  signal W_store_kernel_3131_delayed_1_0_3233_inst_ack_0 : boolean;
  signal phi_stmt_2905_req_0 : boolean;
  signal RPIPE_size_pipe_2883_inst_ack_1 : boolean;
  signal phi_stmt_2905_ack_0 : boolean;
  signal W_store_kernel_3131_delayed_1_0_3233_inst_req_0 : boolean;
  signal n_col_3276_2909_buf_ack_0 : boolean;
  signal nacc1_3293_2894_buf_req_0 : boolean;
  signal nacc1_3293_2894_buf_ack_0 : boolean;
  signal n_col_3276_2909_buf_ack_1 : boolean;
  signal n_col_3276_2909_buf_req_1 : boolean;
  signal SUB_u16_u16_2875_inst_req_0 : boolean;
  signal SUB_u16_u16_3208_inst_ack_0 : boolean;
  signal do_while_stmt_2887_branch_req_0 : boolean;
  signal n_row_3284_2904_buf_req_0 : boolean;
  signal nacc2_3302_2899_buf_ack_0 : boolean;
  signal SUB_u16_u16_2875_inst_ack_0 : boolean;
  signal n_row_3284_2904_buf_ack_1 : boolean;
  signal W_store_kernel_3135_delayed_1_0_3240_inst_req_0 : boolean;
  signal SUB_u16_u16_2885_inst_req_0 : boolean;
  signal W_store_kernel_3127_delayed_1_0_3226_inst_req_1 : boolean;
  signal n_row_3284_2904_buf_ack_0 : boolean;
  signal phi_stmt_2895_req_1 : boolean;
  signal n_row_3284_2904_buf_req_1 : boolean;
  signal W_store_kernel_3127_delayed_1_0_3226_inst_ack_0 : boolean;
  signal phi_stmt_2905_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_3230_inst_req_0 : boolean;
  signal phi_stmt_2900_ack_0 : boolean;
  signal phi_stmt_2900_req_0 : boolean;
  signal phi_stmt_2900_req_1 : boolean;
  signal W_acc2_3079_delayed_1_0_3171_inst_ack_1 : boolean;
  signal nacc2_3302_2899_buf_ack_1 : boolean;
  signal nacc2_3302_2899_buf_req_1 : boolean;
  signal SUB_u16_u16_2885_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_3237_inst_req_1 : boolean;
  signal phi_stmt_2895_req_0 : boolean;
  signal W_acc2_3079_delayed_1_0_3171_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_3237_inst_ack_1 : boolean;
  signal W_acc2_3079_delayed_1_0_3171_inst_ack_0 : boolean;
  signal phi_stmt_2910_req_1 : boolean;
  signal W_read_k_3004_delayed_1_0_3084_inst_ack_0 : boolean;
  signal phi_stmt_2910_req_0 : boolean;
  signal W_acc2_3079_delayed_1_0_3171_inst_req_0 : boolean;
  signal phi_stmt_2910_ack_0 : boolean;
  signal W_acc1_3070_delayed_1_0_3159_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_3237_inst_ack_0 : boolean;
  signal W_acc1_3070_delayed_1_0_3159_inst_req_1 : boolean;
  signal W_acc1_3070_delayed_1_0_3159_inst_ack_0 : boolean;
  signal W_acc1_3070_delayed_1_0_3159_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_3237_inst_req_0 : boolean;
  signal W_read_k_3016_delayed_1_0_3102_inst_ack_1 : boolean;
  signal W_read_k_3016_delayed_1_0_3102_inst_req_1 : boolean;
  signal n_num_3265_2914_buf_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_3230_inst_ack_1 : boolean;
  signal n_num_3265_2914_buf_ack_0 : boolean;
  signal n_num_3265_2914_buf_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_3230_inst_req_1 : boolean;
  signal n_num_3265_2914_buf_ack_1 : boolean;
  signal W_read_k_3016_delayed_1_0_3102_inst_ack_0 : boolean;
  signal W_read_k_3016_delayed_1_0_3102_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_3230_inst_ack_0 : boolean;
  signal phi_stmt_2915_req_1 : boolean;
  signal W_read_k_3010_delayed_1_0_3093_inst_ack_1 : boolean;
  signal W_store_kernel_3131_delayed_1_0_3233_inst_ack_1 : boolean;
  signal phi_stmt_2915_req_0 : boolean;
  signal phi_stmt_2915_ack_0 : boolean;
  signal n_chl_3254_2919_buf_req_0 : boolean;
  signal n_chl_3254_2919_buf_ack_0 : boolean;
  signal n_chl_3254_2919_buf_req_1 : boolean;
  signal n_chl_3254_2919_buf_ack_1 : boolean;
  signal RPIPE_input_pipe1_2932_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_2932_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_2932_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_2932_inst_ack_1 : boolean;
  signal RPIPE_input_pipe2_2936_inst_req_0 : boolean;
  signal RPIPE_input_pipe2_2936_inst_ack_0 : boolean;
  signal RPIPE_input_pipe2_2936_inst_req_1 : boolean;
  signal RPIPE_input_pipe2_2936_inst_ack_1 : boolean;
  signal RPIPE_input_pipe3_2940_inst_req_0 : boolean;
  signal RPIPE_input_pipe3_2940_inst_ack_0 : boolean;
  signal RPIPE_input_pipe3_2940_inst_req_1 : boolean;
  signal RPIPE_input_pipe3_2940_inst_ack_1 : boolean;
  signal RPIPE_input_pipe4_2944_inst_req_0 : boolean;
  signal RPIPE_input_pipe4_2944_inst_ack_0 : boolean;
  signal RPIPE_input_pipe4_2944_inst_req_1 : boolean;
  signal RPIPE_input_pipe4_2944_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2948_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2948_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2948_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2948_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2952_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2952_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2952_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2952_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2956_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2956_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2956_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2956_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2960_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2960_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2960_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2960_inst_ack_1 : boolean;
  signal W_read_ip_2906_delayed_1_0_2962_inst_req_0 : boolean;
  signal W_read_ip_2906_delayed_1_0_2962_inst_ack_0 : boolean;
  signal W_read_ip_2906_delayed_1_0_2962_inst_req_1 : boolean;
  signal W_read_ip_2906_delayed_1_0_2962_inst_ack_1 : boolean;
  signal W_read_ip_2912_delayed_1_0_2971_inst_req_0 : boolean;
  signal W_read_ip_2912_delayed_1_0_2971_inst_ack_0 : boolean;
  signal W_read_ip_2912_delayed_1_0_2971_inst_req_1 : boolean;
  signal W_read_ip_2912_delayed_1_0_2971_inst_ack_1 : boolean;
  signal W_read_ip_2918_delayed_1_0_2980_inst_req_0 : boolean;
  signal W_read_ip_2918_delayed_1_0_2980_inst_ack_0 : boolean;
  signal W_read_ip_2918_delayed_1_0_2980_inst_req_1 : boolean;
  signal W_read_ip_2918_delayed_1_0_2980_inst_ack_1 : boolean;
  signal W_read_ip_2924_delayed_1_0_2989_inst_req_0 : boolean;
  signal W_read_ip_2924_delayed_1_0_2989_inst_ack_0 : boolean;
  signal W_read_ip_2924_delayed_1_0_2989_inst_req_1 : boolean;
  signal W_read_ip_2924_delayed_1_0_2989_inst_ack_1 : boolean;
  signal W_write_input_2938_delayed_1_0_3007_inst_req_0 : boolean;
  signal W_write_input_2938_delayed_1_0_3007_inst_ack_0 : boolean;
  signal W_write_input_2938_delayed_1_0_3007_inst_req_1 : boolean;
  signal W_write_input_2938_delayed_1_0_3007_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_3011_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_3011_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_3011_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_3011_inst_ack_1 : boolean;
  signal W_write_input_2942_delayed_1_0_3014_inst_req_0 : boolean;
  signal W_write_input_2942_delayed_1_0_3014_inst_ack_0 : boolean;
  signal W_write_input_2942_delayed_1_0_3014_inst_req_1 : boolean;
  signal W_write_input_2942_delayed_1_0_3014_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_3018_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_3018_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_3018_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_3018_inst_ack_1 : boolean;
  signal W_write_input_2946_delayed_1_0_3021_inst_req_0 : boolean;
  signal W_write_input_2946_delayed_1_0_3021_inst_ack_0 : boolean;
  signal W_write_input_2946_delayed_1_0_3021_inst_req_1 : boolean;
  signal W_write_input_2946_delayed_1_0_3021_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_3025_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_3025_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_3025_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_3025_inst_ack_1 : boolean;
  signal W_write_input_2950_delayed_1_0_3028_inst_req_0 : boolean;
  signal W_write_input_2950_delayed_1_0_3028_inst_ack_0 : boolean;
  signal W_write_input_2950_delayed_1_0_3028_inst_req_1 : boolean;
  signal W_write_input_2950_delayed_1_0_3028_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_3032_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_3032_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_3032_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_3032_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_3062_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_3062_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_3062_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_3062_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe2_3066_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe2_3066_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_3066_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe2_3066_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe3_3070_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe3_3070_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe3_3070_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe3_3070_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_3074_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_3074_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_3074_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_3074_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_3078_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_3078_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_3078_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_3078_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_3082_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_3082_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_3082_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_3082_inst_ack_1 : boolean;
  signal W_store_kernel_3135_delayed_1_0_3240_inst_ack_0 : boolean;
  signal W_store_kernel_3135_delayed_1_0_3240_inst_req_1 : boolean;
  signal W_store_kernel_3135_delayed_1_0_3240_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_3244_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_3244_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_3244_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_3244_inst_ack_1 : boolean;
  signal W_num_done_3178_delayed_1_0_3285_inst_req_0 : boolean;
  signal W_num_done_3178_delayed_1_0_3285_inst_ack_0 : boolean;
  signal W_num_done_3178_delayed_1_0_3285_inst_req_1 : boolean;
  signal W_num_done_3178_delayed_1_0_3285_inst_ack_1 : boolean;
  signal W_num_done_3184_delayed_1_0_3294_inst_req_0 : boolean;
  signal W_num_done_3184_delayed_1_0_3294_inst_ack_0 : boolean;
  signal W_num_done_3184_delayed_1_0_3294_inst_req_1 : boolean;
  signal W_num_done_3184_delayed_1_0_3294_inst_ack_1 : boolean;
  signal W_num_done_3189_delayed_1_0_3303_inst_req_0 : boolean;
  signal W_num_done_3189_delayed_1_0_3303_inst_ack_0 : boolean;
  signal W_num_done_3189_delayed_1_0_3303_inst_req_1 : boolean;
  signal W_num_done_3189_delayed_1_0_3303_inst_ack_1 : boolean;
  signal type_cast_3309_inst_req_0 : boolean;
  signal type_cast_3309_inst_ack_0 : boolean;
  signal type_cast_3309_inst_req_1 : boolean;
  signal type_cast_3309_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_3307_inst_req_0 : boolean;
  signal WPIPE_output_pipe_3307_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_3307_inst_req_1 : boolean;
  signal WPIPE_output_pipe_3307_inst_ack_1 : boolean;
  signal W_num_done_3194_delayed_1_0_3311_inst_req_0 : boolean;
  signal W_num_done_3194_delayed_1_0_3311_inst_ack_0 : boolean;
  signal W_num_done_3194_delayed_1_0_3311_inst_req_1 : boolean;
  signal W_num_done_3194_delayed_1_0_3311_inst_ack_1 : boolean;
  signal type_cast_3317_inst_req_0 : boolean;
  signal type_cast_3317_inst_ack_0 : boolean;
  signal type_cast_3317_inst_req_1 : boolean;
  signal type_cast_3317_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_3315_inst_req_0 : boolean;
  signal WPIPE_output_pipe_3315_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_3315_inst_req_1 : boolean;
  signal WPIPE_output_pipe_3315_inst_ack_1 : boolean;
  signal do_while_stmt_2887_branch_ack_0 : boolean;
  signal do_while_stmt_2887_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3322_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3322_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_3322_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_3322_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_6745_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_6745_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_6745_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_6745_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_6745: Block -- control-path 
    signal convolve_CP_6745_elements: BooleanArray(323 downto 0);
    -- 
  begin -- 
    convolve_CP_6745_elements(0) <= convolve_CP_6745_start;
    convolve_CP_6745_symbol <= convolve_CP_6745_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	323 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_2870/merge_stmt_2871__entry__
      -- CP-element group 0: 	 branch_block_stmt_2870/branch_block_stmt_2870__entry__
      -- CP-element group 0: 	 branch_block_stmt_2870/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2870/merge_stmt_2871_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_2870/merge_stmt_2871__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_2870/merge_stmt_2871__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_2870/branch_block_stmt_2870__exit__
      -- CP-element group 1: 	 branch_block_stmt_2870/$exit
      -- CP-element group 1: 	 $exit
      -- 
    convolve_CP_6745_elements(1) <= false; 
    -- CP-element group 2:  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	320 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	321 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2870/assign_stmt_3324__entry__
      -- CP-element group 2: 	 branch_block_stmt_2870/do_while_stmt_2887__exit__
      -- CP-element group 2: 	 branch_block_stmt_2870/assign_stmt_3324/$entry
      -- CP-element group 2: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_Sample/req
      -- 
    req_7797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(2), ack => WPIPE_input_done_pipe_3322_inst_req_0); -- 
    convolve_CP_6745_elements(2) <= convolve_CP_6745_elements(320);
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	323 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_sample_completed_
      -- 
    ra_6777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2873_inst_ack_0, ack => convolve_CP_6745_elements(3)); -- 
    cr_6781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(3), ack => RPIPE_num_out_pipe_2873_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_Sample/$entry
      -- 
    ca_6782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2873_inst_ack_1, ack => convolve_CP_6745_elements(4)); -- 
    rr_6804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(4), ack => RPIPE_num_out_pipe_2878_inst_req_0); -- 
    rr_6786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(4), ack => SUB_u16_u16_2875_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_Sample/ra
      -- 
    ra_6787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2875_inst_ack_0, ack => convolve_CP_6745_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	323 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	15 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_update_completed_
      -- 
    ca_6792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2875_inst_ack_1, ack => convolve_CP_6745_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_update_start_
      -- CP-element group 7: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_sample_completed_
      -- 
    ra_6805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2878_inst_ack_0, ack => convolve_CP_6745_elements(7)); -- 
    cr_6809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(7), ack => RPIPE_num_out_pipe_2878_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2878_update_completed_
      -- 
    ca_6810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2878_inst_ack_1, ack => convolve_CP_6745_elements(8)); -- 
    rr_6814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(8), ack => SUB_u16_u16_2880_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_Sample/ra
      -- 
    ra_6815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2880_inst_ack_0, ack => convolve_CP_6745_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	323 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_Update/$exit
      -- 
    ca_6820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2880_inst_ack_1, ack => convolve_CP_6745_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	323 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_update_start_
      -- CP-element group 11: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_Sample/ra
      -- 
    ra_6833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_2883_inst_ack_0, ack => convolve_CP_6745_elements(11)); -- 
    cr_6837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(11), ack => RPIPE_size_pipe_2883_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_Sample/rr
      -- 
    ca_6838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_2883_inst_ack_1, ack => convolve_CP_6745_elements(12)); -- 
    rr_6842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(12), ack => SUB_u16_u16_2885_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_Sample/ra
      -- 
    ra_6843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2885_inst_ack_0, ack => convolve_CP_6745_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	323 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_Update/$exit
      -- 
    ca_6848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2885_inst_ack_1, ack => convolve_CP_6745_elements(14)); -- 
    -- CP-element group 15:  join  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	6 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886__exit__
      -- CP-element group 15: 	 branch_block_stmt_2870/do_while_stmt_2887__entry__
      -- CP-element group 15: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/$exit
      -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(6) & convolve_CP_6745_elements(10) & convolve_CP_6745_elements(14);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887__entry__
      -- CP-element group 16: 	 branch_block_stmt_2870/do_while_stmt_2887/$entry
      -- 
    convolve_CP_6745_elements(16) <= convolve_CP_6745_elements(15);
    -- CP-element group 17:  merge  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	320 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887__exit__
      -- 
    -- Element group convolve_CP_6745_elements(17) is bound as output of CP function.
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2870/do_while_stmt_2887/loop_back
      -- 
    -- Element group convolve_CP_6745_elements(18) is bound as output of CP function.
    -- CP-element group 19:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	318 
    -- CP-element group 19: 	319 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2870/do_while_stmt_2887/condition_done
      -- CP-element group 19: 	 branch_block_stmt_2870/do_while_stmt_2887/loop_exit/$entry
      -- CP-element group 19: 	 branch_block_stmt_2870/do_while_stmt_2887/loop_taken/$entry
      -- 
    convolve_CP_6745_elements(19) <= convolve_CP_6745_elements(24);
    -- CP-element group 20:  branch  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	317 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2870/do_while_stmt_2887/loop_body_done
      -- 
    convolve_CP_6745_elements(20) <= convolve_CP_6745_elements(317);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	109 
    -- CP-element group 21: 	33 
    -- CP-element group 21: 	52 
    -- CP-element group 21: 	90 
    -- CP-element group 21: 	71 
    -- CP-element group 21: 	128 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_6745_elements(21) <= convolve_CP_6745_elements(18);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	35 
    -- CP-element group 22: 	54 
    -- CP-element group 22: 	92 
    -- CP-element group 22: 	73 
    -- CP-element group 22: 	130 
    -- CP-element group 22: 	111 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_6745_elements(22) <= convolve_CP_6745_elements(16);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	65 
    -- CP-element group 23: 	161 
    -- CP-element group 23: 	165 
    -- CP-element group 23: 	149 
    -- CP-element group 23: 	153 
    -- CP-element group 23: 	316 
    -- CP-element group 23: 	29 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	103 
    -- CP-element group 23: 	104 
    -- CP-element group 23: 	122 
    -- CP-element group 23: 	123 
    -- CP-element group 23: 	217 
    -- CP-element group 23: 	221 
    -- CP-element group 23: 	145 
    -- CP-element group 23: 	237 
    -- CP-element group 23: 	261 
    -- CP-element group 23: 	84 
    -- CP-element group 23: 	85 
    -- CP-element group 23: 	66 
    -- CP-element group 23: 	157 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	47 
    -- CP-element group 23: 	141 
    -- CP-element group 23: 	169 
    -- CP-element group 23: 	225 
    -- CP-element group 23: 	229 
    -- CP-element group 23: 	233 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/$entry
      -- CP-element group 23: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_6745_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	316 
    -- CP-element group 24: 	108 
    -- CP-element group 24: 	89 
    -- CP-element group 24: 	70 
    -- CP-element group 24: 	127 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	264 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/condition_evaluated
      -- 
    condition_evaluated_6863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(24), ack => do_while_stmt_2887_branch_req_0); -- 
    convolve_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(316) & convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(127) & convolve_CP_6745_elements(28) & convolve_CP_6745_elements(264);
      gj_convolve_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	65 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	103 
    -- CP-element group 25: 	122 
    -- CP-element group 25: 	84 
    -- CP-element group 25: 	46 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	105 
    -- CP-element group 25: 	124 
    -- CP-element group 25: 	48 
    -- CP-element group 25: 	86 
    -- CP-element group 25: 	67 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/aggregated_phi_sample_req
      -- 
    convolve_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(65) & convolve_CP_6745_elements(29) & convolve_CP_6745_elements(103) & convolve_CP_6745_elements(122) & convolve_CP_6745_elements(84) & convolve_CP_6745_elements(46) & convolve_CP_6745_elements(28);
      gj_convolve_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: 	106 
    -- CP-element group 26: 	125 
    -- CP-element group 26: 	49 
    -- CP-element group 26: 	87 
    -- CP-element group 26: 	68 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	162 
    -- CP-element group 26: 	166 
    -- CP-element group 26: 	150 
    -- CP-element group 26: 	154 
    -- CP-element group 26: 	287 
    -- CP-element group 26: 	291 
    -- CP-element group 26: 	317 
    -- CP-element group 26: 	218 
    -- CP-element group 26: 	222 
    -- CP-element group 26: 	146 
    -- CP-element group 26: 	238 
    -- CP-element group 26: 	242 
    -- CP-element group 26: 	246 
    -- CP-element group 26: 	250 
    -- CP-element group 26: 	254 
    -- CP-element group 26: 	258 
    -- CP-element group 26: 	182 
    -- CP-element group 26: 	186 
    -- CP-element group 26: 	174 
    -- CP-element group 26: 	178 
    -- CP-element group 26: 	158 
    -- CP-element group 26: 	142 
    -- CP-element group 26: 	170 
    -- CP-element group 26: 	226 
    -- CP-element group 26: 	230 
    -- CP-element group 26: 	234 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	65 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	103 
    -- CP-element group 26: 	122 
    -- CP-element group 26: 	84 
    -- CP-element group 26: 	46 
    -- CP-element group 26:  members (7) 
      -- CP-element group 26: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/aggregated_phi_sample_ack
      -- CP-element group 26: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_sample_completed_
      -- 
    convolve_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(31) & convolve_CP_6745_elements(106) & convolve_CP_6745_elements(125) & convolve_CP_6745_elements(49) & convolve_CP_6745_elements(87) & convolve_CP_6745_elements(68);
      gj_convolve_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	104 
    -- CP-element group 27: 	123 
    -- CP-element group 27: 	85 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	47 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	107 
    -- CP-element group 27: 	126 
    -- CP-element group 27: 	50 
    -- CP-element group 27: 	88 
    -- CP-element group 27: 	69 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/aggregated_phi_update_req
      -- 
    convolve_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(30) & convolve_CP_6745_elements(104) & convolve_CP_6745_elements(123) & convolve_CP_6745_elements(85) & convolve_CP_6745_elements(66) & convolve_CP_6745_elements(47);
      gj_convolve_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	32 
    -- CP-element group 28: 	108 
    -- CP-element group 28: 	51 
    -- CP-element group 28: 	89 
    -- CP-element group 28: 	70 
    -- CP-element group 28: 	127 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(32) & convolve_CP_6745_elements(108) & convolve_CP_6745_elements(51) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(127);
      gj_convolve_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	164 
    -- CP-element group 29: 	148 
    -- CP-element group 29: 	152 
    -- CP-element group 29: 	289 
    -- CP-element group 29: 	220 
    -- CP-element group 29: 	144 
    -- CP-element group 29: 	236 
    -- CP-element group 29: 	240 
    -- CP-element group 29: 	244 
    -- CP-element group 29: 	248 
    -- CP-element group 29: 	252 
    -- CP-element group 29: 	256 
    -- CP-element group 29: 	180 
    -- CP-element group 29: 	184 
    -- CP-element group 29: 	176 
    -- CP-element group 29: 	160 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	168 
    -- CP-element group 29: 	224 
    -- CP-element group 29: 	228 
    -- CP-element group 29: 	232 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_sample_start_
      -- 
    convolve_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 1,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(164) & convolve_CP_6745_elements(148) & convolve_CP_6745_elements(152) & convolve_CP_6745_elements(289) & convolve_CP_6745_elements(220) & convolve_CP_6745_elements(144) & convolve_CP_6745_elements(236) & convolve_CP_6745_elements(240) & convolve_CP_6745_elements(244) & convolve_CP_6745_elements(248) & convolve_CP_6745_elements(252) & convolve_CP_6745_elements(256) & convolve_CP_6745_elements(180) & convolve_CP_6745_elements(184) & convolve_CP_6745_elements(176) & convolve_CP_6745_elements(160) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(168) & convolve_CP_6745_elements(224) & convolve_CP_6745_elements(228) & convolve_CP_6745_elements(232);
      gj_convolve_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	255 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	27 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_update_start_
      -- 
    convolve_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(32) & convolve_CP_6745_elements(255);
      gj_convolve_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	26 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_sample_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	253 
    -- CP-element group 32: 	28 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_update_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(32) is bound as output of CP function.
    -- CP-element group 33:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	21 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_loopback_trigger
      -- 
    convolve_CP_6745_elements(33) <= convolve_CP_6745_elements(21);
    -- CP-element group 34:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_loopback_sample_req_ps
      -- CP-element group 34: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_loopback_sample_req
      -- 
    phi_stmt_2889_loopback_sample_req_6878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2889_loopback_sample_req_6878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(34), ack => phi_stmt_2889_req_1); -- 
    -- Element group convolve_CP_6745_elements(34) is bound as output of CP function.
    -- CP-element group 35:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	22 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_entry_trigger
      -- 
    convolve_CP_6745_elements(35) <= convolve_CP_6745_elements(22);
    -- CP-element group 36:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_entry_sample_req_ps
      -- CP-element group 36: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_entry_sample_req
      -- 
    phi_stmt_2889_entry_sample_req_6881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2889_entry_sample_req_6881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(36), ack => phi_stmt_2889_req_0); -- 
    -- Element group convolve_CP_6745_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_phi_mux_ack_ps
      -- CP-element group 37: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2889_phi_mux_ack
      -- 
    phi_stmt_2889_phi_mux_ack_6884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2889_ack_0, ack => convolve_CP_6745_elements(37)); -- 
    -- CP-element group 38:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2893_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2893_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2893_sample_start__ps
      -- CP-element group 38: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2893_sample_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2893_update_start__ps
      -- CP-element group 39: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2893_update_start_
      -- 
    -- Element group convolve_CP_6745_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2893_update_completed__ps
      -- 
    convolve_CP_6745_elements(40) <= convolve_CP_6745_elements(41);
    -- CP-element group 41:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	40 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2893_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => convolve_CP_6745_elements(39), ack => convolve_CP_6745_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_sample_start__ps
      -- CP-element group 42: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_Sample/req
      -- 
    req_6905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(42), ack => nacc1_3293_2894_buf_req_0); -- 
    -- Element group convolve_CP_6745_elements(42) is bound as output of CP function.
    -- CP-element group 43:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_Update/req
      -- CP-element group 43: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_update_start__ps
      -- CP-element group 43: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_update_start_
      -- CP-element group 43: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_Update/$entry
      -- 
    req_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(43), ack => nacc1_3293_2894_buf_req_1); -- 
    -- Element group convolve_CP_6745_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_sample_completed__ps
      -- CP-element group 44: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_Sample/ack
      -- 
    ack_6906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc1_3293_2894_buf_ack_0, ack => convolve_CP_6745_elements(44)); -- 
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_update_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc1_2894_Update/$exit
      -- 
    ack_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc1_3293_2894_buf_ack_1, ack => convolve_CP_6745_elements(45)); -- 
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	164 
    -- CP-element group 46: 	148 
    -- CP-element group 46: 	152 
    -- CP-element group 46: 	293 
    -- CP-element group 46: 	220 
    -- CP-element group 46: 	236 
    -- CP-element group 46: 	240 
    -- CP-element group 46: 	244 
    -- CP-element group 46: 	248 
    -- CP-element group 46: 	252 
    -- CP-element group 46: 	260 
    -- CP-element group 46: 	180 
    -- CP-element group 46: 	184 
    -- CP-element group 46: 	156 
    -- CP-element group 46: 	188 
    -- CP-element group 46: 	26 
    -- CP-element group 46: 	168 
    -- CP-element group 46: 	172 
    -- CP-element group 46: 	224 
    -- CP-element group 46: 	228 
    -- CP-element group 46: 	232 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	25 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_sample_start_
      -- 
    convolve_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(164) & convolve_CP_6745_elements(148) & convolve_CP_6745_elements(152) & convolve_CP_6745_elements(293) & convolve_CP_6745_elements(220) & convolve_CP_6745_elements(236) & convolve_CP_6745_elements(240) & convolve_CP_6745_elements(244) & convolve_CP_6745_elements(248) & convolve_CP_6745_elements(252) & convolve_CP_6745_elements(260) & convolve_CP_6745_elements(180) & convolve_CP_6745_elements(184) & convolve_CP_6745_elements(156) & convolve_CP_6745_elements(188) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(168) & convolve_CP_6745_elements(172) & convolve_CP_6745_elements(224) & convolve_CP_6745_elements(228) & convolve_CP_6745_elements(232);
      gj_convolve_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	23 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	259 
    -- CP-element group 47: 	51 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	27 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_update_start_
      -- 
    convolve_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(259) & convolve_CP_6745_elements(51);
      gj_convolve_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	25 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_sample_start__ps
      -- 
    convolve_CP_6745_elements(48) <= convolve_CP_6745_elements(25);
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	26 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_sample_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	27 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_update_start__ps
      -- 
    convolve_CP_6745_elements(50) <= convolve_CP_6745_elements(27);
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	257 
    -- CP-element group 51: 	28 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	47 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_update_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	21 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_loopback_trigger
      -- 
    convolve_CP_6745_elements(52) <= convolve_CP_6745_elements(21);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_loopback_sample_req
      -- CP-element group 53: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_loopback_sample_req_ps
      -- 
    phi_stmt_2895_loopback_sample_req_6922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2895_loopback_sample_req_6922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(53), ack => phi_stmt_2895_req_1); -- 
    -- Element group convolve_CP_6745_elements(53) is bound as output of CP function.
    -- CP-element group 54:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	22 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_entry_trigger
      -- 
    convolve_CP_6745_elements(54) <= convolve_CP_6745_elements(22);
    -- CP-element group 55:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_entry_sample_req_ps
      -- CP-element group 55: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_entry_sample_req
      -- 
    phi_stmt_2895_entry_sample_req_6925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2895_entry_sample_req_6925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(55), ack => phi_stmt_2895_req_0); -- 
    -- Element group convolve_CP_6745_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_phi_mux_ack_ps
      -- CP-element group 56: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2895_phi_mux_ack
      -- 
    phi_stmt_2895_phi_mux_ack_6928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2895_ack_0, ack => convolve_CP_6745_elements(56)); -- 
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2898_sample_start__ps
      -- CP-element group 57: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2898_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2898_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2898_sample_completed_
      -- 
    -- Element group convolve_CP_6745_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2898_update_start_
      -- CP-element group 58: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2898_update_start__ps
      -- 
    -- Element group convolve_CP_6745_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2898_update_completed__ps
      -- 
    convolve_CP_6745_elements(59) <= convolve_CP_6745_elements(60);
    -- CP-element group 60:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	59 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2898_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => convolve_CP_6745_elements(58), ack => convolve_CP_6745_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_Sample/req
      -- CP-element group 61: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_sample_start__ps
      -- CP-element group 61: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_Sample/$entry
      -- 
    req_6949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(61), ack => nacc2_3302_2899_buf_req_0); -- 
    -- Element group convolve_CP_6745_elements(61) is bound as output of CP function.
    -- CP-element group 62:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_update_start__ps
      -- CP-element group 62: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_Update/req
      -- 
    req_6954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(62), ack => nacc2_3302_2899_buf_req_1); -- 
    -- Element group convolve_CP_6745_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_sample_completed__ps
      -- CP-element group 63: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_Sample/$exit
      -- 
    ack_6950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc2_3302_2899_buf_ack_0, ack => convolve_CP_6745_elements(63)); -- 
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_update_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_nacc2_2899_Update/ack
      -- 
    ack_6955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc2_3302_2899_buf_ack_1, ack => convolve_CP_6745_elements(64)); -- 
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	23 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	26 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	25 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_sample_start_
      -- 
    convolve_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(26);
      gj_convolve_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	23 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	281 
    -- CP-element group 66: 	218 
    -- CP-element group 66: 	222 
    -- CP-element group 66: 	238 
    -- CP-element group 66: 	243 
    -- CP-element group 66: 	247 
    -- CP-element group 66: 	251 
    -- CP-element group 66: 	70 
    -- CP-element group 66: 	226 
    -- CP-element group 66: 	230 
    -- CP-element group 66: 	234 
    -- CP-element group 66: 	267 
    -- CP-element group 66: 	274 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	27 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_update_start_
      -- 
    convolve_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(281) & convolve_CP_6745_elements(218) & convolve_CP_6745_elements(222) & convolve_CP_6745_elements(238) & convolve_CP_6745_elements(243) & convolve_CP_6745_elements(247) & convolve_CP_6745_elements(251) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(226) & convolve_CP_6745_elements(230) & convolve_CP_6745_elements(234) & convolve_CP_6745_elements(267) & convolve_CP_6745_elements(274);
      gj_convolve_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_sample_start__ps
      -- 
    convolve_CP_6745_elements(67) <= convolve_CP_6745_elements(25);
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	26 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_sample_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(68) is bound as output of CP function.
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	27 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_update_start__ps
      -- 
    convolve_CP_6745_elements(69) <= convolve_CP_6745_elements(27);
    -- CP-element group 70:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	218 
    -- CP-element group 70: 	222 
    -- CP-element group 70: 	238 
    -- CP-element group 70: 	241 
    -- CP-element group 70: 	245 
    -- CP-element group 70: 	249 
    -- CP-element group 70: 	24 
    -- CP-element group 70: 	28 
    -- CP-element group 70: 	226 
    -- CP-element group 70: 	230 
    -- CP-element group 70: 	234 
    -- CP-element group 70: 	265 
    -- CP-element group 70: 	272 
    -- CP-element group 70: 	279 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	66 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_update_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(70) is bound as output of CP function.
    -- CP-element group 71:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	21 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_loopback_trigger
      -- 
    convolve_CP_6745_elements(71) <= convolve_CP_6745_elements(21);
    -- CP-element group 72:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_loopback_sample_req_ps
      -- CP-element group 72: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_loopback_sample_req
      -- 
    phi_stmt_2900_loopback_sample_req_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2900_loopback_sample_req_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(72), ack => phi_stmt_2900_req_1); -- 
    -- Element group convolve_CP_6745_elements(72) is bound as output of CP function.
    -- CP-element group 73:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	22 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_entry_trigger
      -- 
    convolve_CP_6745_elements(73) <= convolve_CP_6745_elements(22);
    -- CP-element group 74:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_entry_sample_req_ps
      -- CP-element group 74: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_entry_sample_req
      -- 
    phi_stmt_2900_entry_sample_req_6969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2900_entry_sample_req_6969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(74), ack => phi_stmt_2900_req_0); -- 
    -- Element group convolve_CP_6745_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_phi_mux_ack_ps
      -- CP-element group 75: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2900_phi_mux_ack
      -- 
    phi_stmt_2900_phi_mux_ack_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2900_ack_0, ack => convolve_CP_6745_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2903_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2903_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2903_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2903_sample_start__ps
      -- 
    -- Element group convolve_CP_6745_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2903_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2903_update_start__ps
      -- 
    -- Element group convolve_CP_6745_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2903_update_completed__ps
      -- 
    convolve_CP_6745_elements(78) <= convolve_CP_6745_elements(79);
    -- CP-element group 79:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	78 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2903_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convolve_CP_6745_elements(77), ack => convolve_CP_6745_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_Sample/req
      -- CP-element group 80: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_sample_start__ps
      -- 
    req_6993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(80), ack => n_row_3284_2904_buf_req_0); -- 
    -- Element group convolve_CP_6745_elements(80) is bound as output of CP function.
    -- CP-element group 81:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_update_start_
      -- CP-element group 81: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_update_start__ps
      -- CP-element group 81: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_Update/req
      -- 
    req_6998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(81), ack => n_row_3284_2904_buf_req_1); -- 
    -- Element group convolve_CP_6745_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_sample_completed__ps
      -- CP-element group 82: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_Sample/ack
      -- 
    ack_6994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3284_2904_buf_ack_0, ack => convolve_CP_6745_elements(82)); -- 
    -- CP-element group 83:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_update_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_row_2904_Update/ack
      -- 
    ack_6999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3284_2904_buf_ack_1, ack => convolve_CP_6745_elements(83)); -- 
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	23 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	26 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	25 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_sample_start_
      -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(26);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	23 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	162 
    -- CP-element group 85: 	166 
    -- CP-element group 85: 	150 
    -- CP-element group 85: 	154 
    -- CP-element group 85: 	281 
    -- CP-element group 85: 	218 
    -- CP-element group 85: 	222 
    -- CP-element group 85: 	146 
    -- CP-element group 85: 	238 
    -- CP-element group 85: 	243 
    -- CP-element group 85: 	247 
    -- CP-element group 85: 	251 
    -- CP-element group 85: 	183 
    -- CP-element group 85: 	175 
    -- CP-element group 85: 	179 
    -- CP-element group 85: 	89 
    -- CP-element group 85: 	212 
    -- CP-element group 85: 	158 
    -- CP-element group 85: 	187 
    -- CP-element group 85: 	191 
    -- CP-element group 85: 	142 
    -- CP-element group 85: 	205 
    -- CP-element group 85: 	170 
    -- CP-element group 85: 	198 
    -- CP-element group 85: 	226 
    -- CP-element group 85: 	230 
    -- CP-element group 85: 	234 
    -- CP-element group 85: 	267 
    -- CP-element group 85: 	274 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	27 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_update_start_
      -- 
    convolve_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 29) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_markings: IntegerArray(0 to 29)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_delays: IntegerArray(0 to 29) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 30); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(162) & convolve_CP_6745_elements(166) & convolve_CP_6745_elements(150) & convolve_CP_6745_elements(154) & convolve_CP_6745_elements(281) & convolve_CP_6745_elements(218) & convolve_CP_6745_elements(222) & convolve_CP_6745_elements(146) & convolve_CP_6745_elements(238) & convolve_CP_6745_elements(243) & convolve_CP_6745_elements(247) & convolve_CP_6745_elements(251) & convolve_CP_6745_elements(183) & convolve_CP_6745_elements(175) & convolve_CP_6745_elements(179) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(212) & convolve_CP_6745_elements(158) & convolve_CP_6745_elements(187) & convolve_CP_6745_elements(191) & convolve_CP_6745_elements(142) & convolve_CP_6745_elements(205) & convolve_CP_6745_elements(170) & convolve_CP_6745_elements(198) & convolve_CP_6745_elements(226) & convolve_CP_6745_elements(230) & convolve_CP_6745_elements(234) & convolve_CP_6745_elements(267) & convolve_CP_6745_elements(274);
      gj_convolve_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 30, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	25 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_sample_start__ps
      -- 
    convolve_CP_6745_elements(86) <= convolve_CP_6745_elements(25);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	26 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_sample_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(87) is bound as output of CP function.
    -- CP-element group 88:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	27 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_update_start__ps
      -- 
    convolve_CP_6745_elements(88) <= convolve_CP_6745_elements(27);
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	162 
    -- CP-element group 89: 	166 
    -- CP-element group 89: 	150 
    -- CP-element group 89: 	154 
    -- CP-element group 89: 	218 
    -- CP-element group 89: 	222 
    -- CP-element group 89: 	146 
    -- CP-element group 89: 	238 
    -- CP-element group 89: 	241 
    -- CP-element group 89: 	245 
    -- CP-element group 89: 	249 
    -- CP-element group 89: 	181 
    -- CP-element group 89: 	185 
    -- CP-element group 89: 	177 
    -- CP-element group 89: 	158 
    -- CP-element group 89: 	189 
    -- CP-element group 89: 	203 
    -- CP-element group 89: 	24 
    -- CP-element group 89: 	28 
    -- CP-element group 89: 	142 
    -- CP-element group 89: 	210 
    -- CP-element group 89: 	170 
    -- CP-element group 89: 	173 
    -- CP-element group 89: 	196 
    -- CP-element group 89: 	226 
    -- CP-element group 89: 	230 
    -- CP-element group 89: 	234 
    -- CP-element group 89: 	265 
    -- CP-element group 89: 	272 
    -- CP-element group 89: 	279 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	85 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_update_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(89) is bound as output of CP function.
    -- CP-element group 90:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	21 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_loopback_trigger
      -- 
    convolve_CP_6745_elements(90) <= convolve_CP_6745_elements(21);
    -- CP-element group 91:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_loopback_sample_req_ps
      -- CP-element group 91: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_loopback_sample_req
      -- 
    phi_stmt_2905_loopback_sample_req_7010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2905_loopback_sample_req_7010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(91), ack => phi_stmt_2905_req_1); -- 
    -- Element group convolve_CP_6745_elements(91) is bound as output of CP function.
    -- CP-element group 92:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	22 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_entry_trigger
      -- 
    convolve_CP_6745_elements(92) <= convolve_CP_6745_elements(22);
    -- CP-element group 93:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_entry_sample_req
      -- CP-element group 93: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_entry_sample_req_ps
      -- 
    phi_stmt_2905_entry_sample_req_7013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2905_entry_sample_req_7013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(93), ack => phi_stmt_2905_req_0); -- 
    -- Element group convolve_CP_6745_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_phi_mux_ack
      -- CP-element group 94: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2905_phi_mux_ack_ps
      -- 
    phi_stmt_2905_phi_mux_ack_7016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2905_ack_0, ack => convolve_CP_6745_elements(94)); -- 
    -- CP-element group 95:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2908_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2908_sample_start__ps
      -- CP-element group 95: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2908_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2908_sample_start_
      -- 
    -- Element group convolve_CP_6745_elements(95) is bound as output of CP function.
    -- CP-element group 96:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2908_update_start__ps
      -- CP-element group 96: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2908_update_start_
      -- 
    -- Element group convolve_CP_6745_elements(96) is bound as output of CP function.
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2908_update_completed__ps
      -- 
    convolve_CP_6745_elements(97) <= convolve_CP_6745_elements(98);
    -- CP-element group 98:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	97 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2908_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(98) is a control-delay.
    cp_element_98_delay: control_delay_element  generic map(name => " 98_delay", delay_value => 1)  port map(req => convolve_CP_6745_elements(96), ack => convolve_CP_6745_elements(98), clk => clk, reset =>reset);
    -- CP-element group 99:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (4) 
      -- CP-element group 99: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_sample_start__ps
      -- CP-element group 99: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_Sample/req
      -- CP-element group 99: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_Sample/$entry
      -- 
    req_7037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(99), ack => n_col_3276_2909_buf_req_0); -- 
    -- Element group convolve_CP_6745_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_update_start__ps
      -- CP-element group 100: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_Update/$entry
      -- 
    req_7042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(100), ack => n_col_3276_2909_buf_req_1); -- 
    -- Element group convolve_CP_6745_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_sample_completed__ps
      -- CP-element group 101: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_Sample/ack
      -- CP-element group 101: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_sample_completed_
      -- 
    ack_7038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3276_2909_buf_ack_0, ack => convolve_CP_6745_elements(101)); -- 
    -- CP-element group 102:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_update_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_Update/ack
      -- CP-element group 102: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_col_2909_Update/$exit
      -- 
    ack_7043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3276_2909_buf_ack_1, ack => convolve_CP_6745_elements(102)); -- 
    -- CP-element group 103:  join  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	23 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	26 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	25 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_sample_start_
      -- 
    convolve_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(26);
      gj_convolve_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	23 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	162 
    -- CP-element group 104: 	166 
    -- CP-element group 104: 	150 
    -- CP-element group 104: 	154 
    -- CP-element group 104: 	288 
    -- CP-element group 104: 	292 
    -- CP-element group 104: 	296 
    -- CP-element group 104: 	307 
    -- CP-element group 104: 	108 
    -- CP-element group 104: 	146 
    -- CP-element group 104: 	183 
    -- CP-element group 104: 	175 
    -- CP-element group 104: 	179 
    -- CP-element group 104: 	212 
    -- CP-element group 104: 	158 
    -- CP-element group 104: 	187 
    -- CP-element group 104: 	191 
    -- CP-element group 104: 	142 
    -- CP-element group 104: 	205 
    -- CP-element group 104: 	170 
    -- CP-element group 104: 	198 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	27 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_update_start_
      -- 
    convolve_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(162) & convolve_CP_6745_elements(166) & convolve_CP_6745_elements(150) & convolve_CP_6745_elements(154) & convolve_CP_6745_elements(288) & convolve_CP_6745_elements(292) & convolve_CP_6745_elements(296) & convolve_CP_6745_elements(307) & convolve_CP_6745_elements(108) & convolve_CP_6745_elements(146) & convolve_CP_6745_elements(183) & convolve_CP_6745_elements(175) & convolve_CP_6745_elements(179) & convolve_CP_6745_elements(212) & convolve_CP_6745_elements(158) & convolve_CP_6745_elements(187) & convolve_CP_6745_elements(191) & convolve_CP_6745_elements(142) & convolve_CP_6745_elements(205) & convolve_CP_6745_elements(170) & convolve_CP_6745_elements(198);
      gj_convolve_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	25 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_sample_start__ps
      -- 
    convolve_CP_6745_elements(105) <= convolve_CP_6745_elements(25);
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	26 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_sample_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(106) is bound as output of CP function.
    -- CP-element group 107:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	27 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_update_start__ps
      -- 
    convolve_CP_6745_elements(107) <= convolve_CP_6745_elements(27);
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	162 
    -- CP-element group 108: 	166 
    -- CP-element group 108: 	150 
    -- CP-element group 108: 	154 
    -- CP-element group 108: 	286 
    -- CP-element group 108: 	290 
    -- CP-element group 108: 	294 
    -- CP-element group 108: 	305 
    -- CP-element group 108: 	146 
    -- CP-element group 108: 	181 
    -- CP-element group 108: 	185 
    -- CP-element group 108: 	177 
    -- CP-element group 108: 	158 
    -- CP-element group 108: 	189 
    -- CP-element group 108: 	203 
    -- CP-element group 108: 	24 
    -- CP-element group 108: 	28 
    -- CP-element group 108: 	142 
    -- CP-element group 108: 	210 
    -- CP-element group 108: 	170 
    -- CP-element group 108: 	173 
    -- CP-element group 108: 	196 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	104 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_update_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(108) is bound as output of CP function.
    -- CP-element group 109:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	21 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_loopback_trigger
      -- 
    convolve_CP_6745_elements(109) <= convolve_CP_6745_elements(21);
    -- CP-element group 110:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_loopback_sample_req
      -- CP-element group 110: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_loopback_sample_req_ps
      -- 
    phi_stmt_2910_loopback_sample_req_7054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2910_loopback_sample_req_7054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(110), ack => phi_stmt_2910_req_1); -- 
    -- Element group convolve_CP_6745_elements(110) is bound as output of CP function.
    -- CP-element group 111:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	22 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_entry_trigger
      -- 
    convolve_CP_6745_elements(111) <= convolve_CP_6745_elements(22);
    -- CP-element group 112:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_entry_sample_req
      -- CP-element group 112: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_entry_sample_req_ps
      -- 
    phi_stmt_2910_entry_sample_req_7057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2910_entry_sample_req_7057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(112), ack => phi_stmt_2910_req_0); -- 
    -- Element group convolve_CP_6745_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_phi_mux_ack
      -- CP-element group 113: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2910_phi_mux_ack_ps
      -- 
    phi_stmt_2910_phi_mux_ack_7060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2910_ack_0, ack => convolve_CP_6745_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2913_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2913_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2913_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2913_sample_completed_
      -- 
    -- Element group convolve_CP_6745_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2913_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2913_update_start_
      -- 
    -- Element group convolve_CP_6745_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2913_update_completed__ps
      -- 
    convolve_CP_6745_elements(116) <= convolve_CP_6745_elements(117);
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2913_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => convolve_CP_6745_elements(115), ack => convolve_CP_6745_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_sample_start__ps
      -- CP-element group 118: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_Sample/req
      -- 
    req_7081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(118), ack => n_num_3265_2914_buf_req_0); -- 
    -- Element group convolve_CP_6745_elements(118) is bound as output of CP function.
    -- CP-element group 119:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_update_start__ps
      -- CP-element group 119: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_update_start_
      -- CP-element group 119: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_Update/req
      -- 
    req_7086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(119), ack => n_num_3265_2914_buf_req_1); -- 
    -- Element group convolve_CP_6745_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (4) 
      -- CP-element group 120: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_sample_completed__ps
      -- CP-element group 120: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_Sample/ack
      -- 
    ack_7082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_3265_2914_buf_ack_0, ack => convolve_CP_6745_elements(120)); -- 
    -- CP-element group 121:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_num_2914_Update/ack
      -- 
    ack_7087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_3265_2914_buf_ack_1, ack => convolve_CP_6745_elements(121)); -- 
    -- CP-element group 122:  join  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	23 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	26 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	25 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_sample_start_
      -- 
    convolve_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(26);
      gj_convolve_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	23 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	288 
    -- CP-element group 123: 	292 
    -- CP-element group 123: 	296 
    -- CP-element group 123: 	307 
    -- CP-element group 123: 	127 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	27 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_update_start_
      -- 
    convolve_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(288) & convolve_CP_6745_elements(292) & convolve_CP_6745_elements(296) & convolve_CP_6745_elements(307) & convolve_CP_6745_elements(127);
      gj_convolve_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	25 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_sample_start__ps
      -- 
    convolve_CP_6745_elements(124) <= convolve_CP_6745_elements(25);
    -- CP-element group 125:  join  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	26 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_sample_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	27 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_update_start__ps
      -- 
    convolve_CP_6745_elements(126) <= convolve_CP_6745_elements(27);
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	286 
    -- CP-element group 127: 	290 
    -- CP-element group 127: 	294 
    -- CP-element group 127: 	305 
    -- CP-element group 127: 	24 
    -- CP-element group 127: 	28 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	123 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_update_completed__ps
      -- 
    -- Element group convolve_CP_6745_elements(127) is bound as output of CP function.
    -- CP-element group 128:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	21 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_loopback_trigger
      -- 
    convolve_CP_6745_elements(128) <= convolve_CP_6745_elements(21);
    -- CP-element group 129:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_loopback_sample_req
      -- CP-element group 129: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_loopback_sample_req_ps
      -- 
    phi_stmt_2915_loopback_sample_req_7098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2915_loopback_sample_req_7098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(129), ack => phi_stmt_2915_req_1); -- 
    -- Element group convolve_CP_6745_elements(129) is bound as output of CP function.
    -- CP-element group 130:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	22 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_entry_trigger
      -- 
    convolve_CP_6745_elements(130) <= convolve_CP_6745_elements(22);
    -- CP-element group 131:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_entry_sample_req
      -- CP-element group 131: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_entry_sample_req_ps
      -- 
    phi_stmt_2915_entry_sample_req_7101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2915_entry_sample_req_7101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(131), ack => phi_stmt_2915_req_0); -- 
    -- Element group convolve_CP_6745_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_phi_mux_ack
      -- CP-element group 132: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/phi_stmt_2915_phi_mux_ack_ps
      -- 
    phi_stmt_2915_phi_mux_ack_7104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2915_ack_0, ack => convolve_CP_6745_elements(132)); -- 
    -- CP-element group 133:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2918_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2918_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2918_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2918_sample_completed_
      -- 
    -- Element group convolve_CP_6745_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2918_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2918_update_start_
      -- 
    -- Element group convolve_CP_6745_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2918_update_completed__ps
      -- 
    convolve_CP_6745_elements(135) <= convolve_CP_6745_elements(136);
    -- CP-element group 136:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	135 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_2918_update_completed_
      -- 
    -- Element group convolve_CP_6745_elements(136) is a control-delay.
    cp_element_136_delay: control_delay_element  generic map(name => " 136_delay", delay_value => 1)  port map(req => convolve_CP_6745_elements(134), ack => convolve_CP_6745_elements(136), clk => clk, reset =>reset);
    -- CP-element group 137:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_sample_start__ps
      -- CP-element group 137: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_Sample/req
      -- 
    req_7125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(137), ack => n_chl_3254_2919_buf_req_0); -- 
    -- Element group convolve_CP_6745_elements(137) is bound as output of CP function.
    -- CP-element group 138:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_update_start__ps
      -- CP-element group 138: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_update_start_
      -- CP-element group 138: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_Update/req
      -- 
    req_7130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(138), ack => n_chl_3254_2919_buf_req_1); -- 
    -- Element group convolve_CP_6745_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_sample_completed__ps
      -- CP-element group 139: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_Sample/ack
      -- 
    ack_7126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3254_2919_buf_ack_0, ack => convolve_CP_6745_elements(139)); -- 
    -- CP-element group 140:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_update_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/R_n_chl_2919_Update/ack
      -- 
    ack_7131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3254_2919_buf_ack_1, ack => convolve_CP_6745_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	23 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	144 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_Sample/rr
      -- 
    rr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(141), ack => RPIPE_input_pipe1_2932_inst_req_0); -- 
    convolve_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(144);
      gj_convolve_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	108 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	89 
    -- CP-element group 142: 	26 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	300 
    -- CP-element group 142: 	194 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	104 
    -- CP-element group 142: 	85 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_update_start_
      -- CP-element group 142: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_Update/cr
      -- 
    cr_7145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(142), ack => RPIPE_input_pipe1_2932_inst_req_1); -- 
    convolve_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 15,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(143) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(194);
      gj_convolve_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_Sample/ra
      -- 
    ra_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_2932_inst_ack_0, ack => convolve_CP_6745_elements(143)); -- 
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	298 
    -- CP-element group 144: 	193 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	29 
    -- CP-element group 144: 	141 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe1_2932_Update/ca
      -- 
    ca_7146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_2932_inst_ack_1, ack => convolve_CP_6745_elements(144)); -- 
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	23 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	148 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_Sample/rr
      -- 
    rr_7154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(145), ack => RPIPE_input_pipe2_2936_inst_req_0); -- 
    convolve_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(148);
      gj_convolve_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	108 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	89 
    -- CP-element group 146: 	26 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	300 
    -- CP-element group 146: 	311 
    -- CP-element group 146: 	201 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	104 
    -- CP-element group 146: 	85 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_update_start_
      -- CP-element group 146: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_Update/cr
      -- 
    cr_7159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(146), ack => RPIPE_input_pipe2_2936_inst_req_1); -- 
    convolve_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(147) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(201);
      gj_convolve_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_Sample/ra
      -- 
    ra_7155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_2936_inst_ack_0, ack => convolve_CP_6745_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	298 
    -- CP-element group 148: 	309 
    -- CP-element group 148: 	200 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	29 
    -- CP-element group 148: 	145 
    -- CP-element group 148: 	46 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe2_2936_Update/ca
      -- 
    ca_7160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_2936_inst_ack_1, ack => convolve_CP_6745_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	23 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	152 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_Sample/rr
      -- 
    rr_7168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(149), ack => RPIPE_input_pipe3_2940_inst_req_0); -- 
    convolve_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(152);
      gj_convolve_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	108 
    -- CP-element group 150: 	89 
    -- CP-element group 150: 	26 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	300 
    -- CP-element group 150: 	311 
    -- CP-element group 150: 	208 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	104 
    -- CP-element group 150: 	85 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_update_start_
      -- CP-element group 150: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_Update/cr
      -- 
    cr_7173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(150), ack => RPIPE_input_pipe3_2940_inst_req_1); -- 
    convolve_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(151) & convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(208);
      gj_convolve_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	150 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_Sample/ra
      -- 
    ra_7169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_2940_inst_ack_0, ack => convolve_CP_6745_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	298 
    -- CP-element group 152: 	309 
    -- CP-element group 152: 	207 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	149 
    -- CP-element group 152: 	29 
    -- CP-element group 152: 	46 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe3_2940_Update/ca
      -- 
    ca_7174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_2940_inst_ack_1, ack => convolve_CP_6745_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	23 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	156 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_Sample/rr
      -- 
    rr_7182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(153), ack => RPIPE_input_pipe4_2944_inst_req_0); -- 
    convolve_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(156);
      gj_convolve_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	108 
    -- CP-element group 154: 	89 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	26 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	311 
    -- CP-element group 154: 	215 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	104 
    -- CP-element group 154: 	85 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_update_start_
      -- CP-element group 154: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_Update/cr
      -- 
    cr_7187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(154), ack => RPIPE_input_pipe4_2944_inst_req_1); -- 
    convolve_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(155) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(215);
      gj_convolve_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	154 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_Sample/ra
      -- 
    ra_7183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe4_2944_inst_ack_0, ack => convolve_CP_6745_elements(155)); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	309 
    -- CP-element group 156: 	214 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	153 
    -- CP-element group 156: 	46 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_input_pipe4_2944_Update/ca
      -- 
    ca_7188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe4_2944_inst_ack_1, ack => convolve_CP_6745_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	23 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	160 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_Sample/rr
      -- 
    rr_7196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(157), ack => RPIPE_xxconvolvexxconv_ip1_2948_inst_req_0); -- 
    convolve_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(160);
      gj_convolve_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	108 
    -- CP-element group 158: 	89 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	26 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	300 
    -- CP-element group 158: 	194 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	104 
    -- CP-element group 158: 	85 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_update_start_
      -- CP-element group 158: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_Update/cr
      -- 
    cr_7201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(158), ack => RPIPE_xxconvolvexxconv_ip1_2948_inst_req_1); -- 
    convolve_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(159) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(194);
      gj_convolve_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	158 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_Sample/ra
      -- 
    ra_7197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_2948_inst_ack_0, ack => convolve_CP_6745_elements(159)); -- 
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	298 
    -- CP-element group 160: 	193 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	29 
    -- CP-element group 160: 	157 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip1_2948_Update/ca
      -- 
    ca_7202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_2948_inst_ack_1, ack => convolve_CP_6745_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	23 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	164 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_Sample/rr
      -- 
    rr_7210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(161), ack => RPIPE_xxconvolvexxconv_ip2_2952_inst_req_0); -- 
    convolve_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(164);
      gj_convolve_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	108 
    -- CP-element group 162: 	89 
    -- CP-element group 162: 	26 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	300 
    -- CP-element group 162: 	311 
    -- CP-element group 162: 	201 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	104 
    -- CP-element group 162: 	85 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_update_start_
      -- CP-element group 162: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_Update/cr
      -- 
    cr_7215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(162), ack => RPIPE_xxconvolvexxconv_ip2_2952_inst_req_1); -- 
    convolve_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(163) & convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(201);
      gj_convolve_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	162 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_Sample/ra
      -- 
    ra_7211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_2952_inst_ack_0, ack => convolve_CP_6745_elements(163)); -- 
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	298 
    -- CP-element group 164: 	309 
    -- CP-element group 164: 	200 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	161 
    -- CP-element group 164: 	29 
    -- CP-element group 164: 	46 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip2_2952_Update/ca
      -- 
    ca_7216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_2952_inst_ack_1, ack => convolve_CP_6745_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	23 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	168 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_Sample/rr
      -- 
    rr_7224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(165), ack => RPIPE_xxconvolvexxconv_ip3_2956_inst_req_0); -- 
    convolve_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(168);
      gj_convolve_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	108 
    -- CP-element group 166: 	89 
    -- CP-element group 166: 	26 
    -- CP-element group 166: 	167 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	300 
    -- CP-element group 166: 	311 
    -- CP-element group 166: 	208 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	104 
    -- CP-element group 166: 	85 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_update_start_
      -- CP-element group 166: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_Update/cr
      -- 
    cr_7229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(166), ack => RPIPE_xxconvolvexxconv_ip3_2956_inst_req_1); -- 
    convolve_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(167) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(208);
      gj_convolve_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	166 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_Sample/ra
      -- 
    ra_7225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_2956_inst_ack_0, ack => convolve_CP_6745_elements(167)); -- 
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	298 
    -- CP-element group 168: 	309 
    -- CP-element group 168: 	207 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	165 
    -- CP-element group 168: 	29 
    -- CP-element group 168: 	46 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip3_2956_Update/ca
      -- 
    ca_7230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_2956_inst_ack_1, ack => convolve_CP_6745_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	23 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	172 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_Sample/rr
      -- 
    rr_7238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(169), ack => RPIPE_xxconvolvexxconv_ip4_2960_inst_req_0); -- 
    convolve_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(172);
      gj_convolve_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	108 
    -- CP-element group 170: 	89 
    -- CP-element group 170: 	26 
    -- CP-element group 170: 	171 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	311 
    -- CP-element group 170: 	215 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	104 
    -- CP-element group 170: 	85 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_update_start_
      -- CP-element group 170: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_Update/cr
      -- 
    cr_7243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(170), ack => RPIPE_xxconvolvexxconv_ip4_2960_inst_req_1); -- 
    convolve_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(171) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(215);
      gj_convolve_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	170 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_Sample/ra
      -- 
    ra_7239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip4_2960_inst_ack_0, ack => convolve_CP_6745_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	309 
    -- CP-element group 172: 	214 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	46 
    -- CP-element group 172: 	169 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_ip4_2960_Update/ca
      -- 
    ca_7244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip4_2960_inst_ack_1, ack => convolve_CP_6745_elements(172)); -- 
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	108 
    -- CP-element group 173: 	89 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_Sample/req
      -- 
    req_7252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(173), ack => W_read_ip_2906_delayed_1_0_2962_inst_req_0); -- 
    convolve_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(175);
      gj_convolve_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	26 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	300 
    -- CP-element group 174: 	176 
    -- CP-element group 174: 	194 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_update_start_
      -- CP-element group 174: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_Update/req
      -- 
    req_7257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(174), ack => W_read_ip_2906_delayed_1_0_2962_inst_req_1); -- 
    convolve_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(176) & convolve_CP_6745_elements(194);
      gj_convolve_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	104 
    -- CP-element group 175: 	85 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_Sample/ack
      -- 
    ack_7253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2906_delayed_1_0_2962_inst_ack_0, ack => convolve_CP_6745_elements(175)); -- 
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	298 
    -- CP-element group 176: 	193 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	29 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2964_Update/ack
      -- 
    ack_7258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2906_delayed_1_0_2962_inst_ack_1, ack => convolve_CP_6745_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	108 
    -- CP-element group 177: 	89 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_Sample/req
      -- 
    req_7266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(177), ack => W_read_ip_2912_delayed_1_0_2971_inst_req_0); -- 
    convolve_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(179);
      gj_convolve_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	26 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	300 
    -- CP-element group 178: 	311 
    -- CP-element group 178: 	180 
    -- CP-element group 178: 	201 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_update_start_
      -- CP-element group 178: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_Update/req
      -- 
    req_7271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(178), ack => W_read_ip_2912_delayed_1_0_2971_inst_req_1); -- 
    convolve_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(180) & convolve_CP_6745_elements(201);
      gj_convolve_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	104 
    -- CP-element group 179: 	177 
    -- CP-element group 179: 	85 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_Sample/ack
      -- 
    ack_7267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2912_delayed_1_0_2971_inst_ack_0, ack => convolve_CP_6745_elements(179)); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	298 
    -- CP-element group 180: 	309 
    -- CP-element group 180: 	200 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	29 
    -- CP-element group 180: 	178 
    -- CP-element group 180: 	46 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2973_Update/ack
      -- 
    ack_7272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2912_delayed_1_0_2971_inst_ack_1, ack => convolve_CP_6745_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	108 
    -- CP-element group 181: 	89 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_Sample/req
      -- 
    req_7280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(181), ack => W_read_ip_2918_delayed_1_0_2980_inst_req_0); -- 
    convolve_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(183);
      gj_convolve_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	26 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	300 
    -- CP-element group 182: 	311 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	208 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_update_start_
      -- CP-element group 182: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_Update/req
      -- 
    req_7285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(182), ack => W_read_ip_2918_delayed_1_0_2980_inst_req_1); -- 
    convolve_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(184) & convolve_CP_6745_elements(208);
      gj_convolve_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	104 
    -- CP-element group 183: 	181 
    -- CP-element group 183: 	85 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_Sample/ack
      -- 
    ack_7281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2918_delayed_1_0_2980_inst_ack_0, ack => convolve_CP_6745_elements(183)); -- 
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	298 
    -- CP-element group 184: 	309 
    -- CP-element group 184: 	207 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	29 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	46 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2982_Update/ack
      -- 
    ack_7286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2918_delayed_1_0_2980_inst_ack_1, ack => convolve_CP_6745_elements(184)); -- 
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	108 
    -- CP-element group 185: 	89 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_Sample/req
      -- 
    req_7294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(185), ack => W_read_ip_2924_delayed_1_0_2989_inst_req_0); -- 
    convolve_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(187);
      gj_convolve_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	26 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	311 
    -- CP-element group 186: 	215 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_update_start_
      -- CP-element group 186: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_Update/req
      -- 
    req_7299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(186), ack => W_read_ip_2924_delayed_1_0_2989_inst_req_1); -- 
    convolve_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(215) & convolve_CP_6745_elements(188);
      gj_convolve_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	104 
    -- CP-element group 187: 	185 
    -- CP-element group 187: 	85 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_Sample/ack
      -- 
    ack_7295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2924_delayed_1_0_2989_inst_ack_0, ack => convolve_CP_6745_elements(187)); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	309 
    -- CP-element group 188: 	214 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: 	46 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_2991_Update/ack
      -- 
    ack_7300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2924_delayed_1_0_2989_inst_ack_1, ack => convolve_CP_6745_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	108 
    -- CP-element group 189: 	89 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_Sample/req
      -- 
    req_7308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(189), ack => W_write_input_2938_delayed_1_0_3007_inst_req_0); -- 
    convolve_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(191);
      gj_convolve_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_update_start_
      -- CP-element group 190: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_Update/req
      -- 
    req_7313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(190), ack => W_write_input_2938_delayed_1_0_3007_inst_req_1); -- 
    convolve_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(192) & convolve_CP_6745_elements(194);
      gj_convolve_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	104 
    -- CP-element group 191: 	85 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_Sample/ack
      -- 
    ack_7309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2938_delayed_1_0_3007_inst_ack_0, ack => convolve_CP_6745_elements(191)); -- 
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3009_Update/ack
      -- 
    ack_7314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2938_delayed_1_0_3007_inst_ack_1, ack => convolve_CP_6745_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	144 
    -- CP-element group 193: 	176 
    -- CP-element group 193: 	160 
    -- CP-element group 193: 	192 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_Sample/req
      -- 
    req_7322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(193), ack => WPIPE_xxconvolvexxconv_ip1_3011_inst_req_0); -- 
    convolve_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(144) & convolve_CP_6745_elements(176) & convolve_CP_6745_elements(160) & convolve_CP_6745_elements(192) & convolve_CP_6745_elements(195);
      gj_convolve_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	174 
    -- CP-element group 194: 	158 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	142 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_update_start_
      -- CP-element group 194: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_Update/req
      -- 
    ack_7323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_3011_inst_ack_0, ack => convolve_CP_6745_elements(194)); -- 
    req_7327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(194), ack => WPIPE_xxconvolvexxconv_ip1_3011_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	317 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip1_3011_Update/ack
      -- 
    ack_7328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_3011_inst_ack_1, ack => convolve_CP_6745_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	108 
    -- CP-element group 196: 	89 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_Sample/req
      -- 
    req_7336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(196), ack => W_write_input_2942_delayed_1_0_3014_inst_req_0); -- 
    convolve_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(198);
      gj_convolve_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_update_start_
      -- CP-element group 197: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_Update/req
      -- 
    req_7341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(197), ack => W_write_input_2942_delayed_1_0_3014_inst_req_1); -- 
    convolve_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(199) & convolve_CP_6745_elements(201);
      gj_convolve_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	104 
    -- CP-element group 198: 	85 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_Sample/ack
      -- 
    ack_7337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2942_delayed_1_0_3014_inst_ack_0, ack => convolve_CP_6745_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3016_Update/ack
      -- 
    ack_7342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2942_delayed_1_0_3014_inst_ack_1, ack => convolve_CP_6745_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	164 
    -- CP-element group 200: 	148 
    -- CP-element group 200: 	180 
    -- CP-element group 200: 	199 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_Sample/req
      -- 
    req_7350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(200), ack => WPIPE_xxconvolvexxconv_ip2_3018_inst_req_0); -- 
    convolve_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(164) & convolve_CP_6745_elements(148) & convolve_CP_6745_elements(180) & convolve_CP_6745_elements(199) & convolve_CP_6745_elements(202);
      gj_convolve_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	162 
    -- CP-element group 201: 	146 
    -- CP-element group 201: 	178 
    -- CP-element group 201: 	197 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_update_start_
      -- CP-element group 201: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_Update/req
      -- 
    ack_7351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_3018_inst_ack_0, ack => convolve_CP_6745_elements(201)); -- 
    req_7355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(201), ack => WPIPE_xxconvolvexxconv_ip2_3018_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	317 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip2_3018_Update/ack
      -- 
    ack_7356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_3018_inst_ack_1, ack => convolve_CP_6745_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	108 
    -- CP-element group 203: 	89 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_Sample/req
      -- 
    req_7364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(203), ack => W_write_input_2946_delayed_1_0_3021_inst_req_0); -- 
    convolve_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(205);
      gj_convolve_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: 	208 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_update_start_
      -- CP-element group 204: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_Update/req
      -- 
    req_7369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(204), ack => W_write_input_2946_delayed_1_0_3021_inst_req_1); -- 
    convolve_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(206) & convolve_CP_6745_elements(208);
      gj_convolve_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	104 
    -- CP-element group 205: 	85 
    -- CP-element group 205: 	203 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_Sample/ack
      -- 
    ack_7365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2946_delayed_1_0_3021_inst_ack_0, ack => convolve_CP_6745_elements(205)); -- 
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3023_Update/ack
      -- 
    ack_7370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2946_delayed_1_0_3021_inst_ack_1, ack => convolve_CP_6745_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	152 
    -- CP-element group 207: 	184 
    -- CP-element group 207: 	206 
    -- CP-element group 207: 	168 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_Sample/req
      -- 
    req_7378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(207), ack => WPIPE_xxconvolvexxconv_ip3_3025_inst_req_0); -- 
    convolve_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(152) & convolve_CP_6745_elements(184) & convolve_CP_6745_elements(206) & convolve_CP_6745_elements(168) & convolve_CP_6745_elements(209);
      gj_convolve_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	166 
    -- CP-element group 208: 	150 
    -- CP-element group 208: 	182 
    -- CP-element group 208: 	204 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_update_start_
      -- CP-element group 208: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_Sample/ack
      -- CP-element group 208: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_Update/req
      -- 
    ack_7379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_3025_inst_ack_0, ack => convolve_CP_6745_elements(208)); -- 
    req_7383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(208), ack => WPIPE_xxconvolvexxconv_ip3_3025_inst_req_1); -- 
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	317 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip3_3025_Update/ack
      -- 
    ack_7384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_3025_inst_ack_1, ack => convolve_CP_6745_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	108 
    -- CP-element group 210: 	89 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_Sample/req
      -- 
    req_7392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(210), ack => W_write_input_2950_delayed_1_0_3028_inst_req_0); -- 
    convolve_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(212);
      gj_convolve_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: 	215 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_update_start_
      -- CP-element group 211: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_Update/req
      -- 
    req_7397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(211), ack => W_write_input_2950_delayed_1_0_3028_inst_req_1); -- 
    convolve_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(213) & convolve_CP_6745_elements(215);
      gj_convolve_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	104 
    -- CP-element group 212: 	85 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_Sample/ack
      -- 
    ack_7393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2950_delayed_1_0_3028_inst_ack_0, ack => convolve_CP_6745_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3030_Update/ack
      -- 
    ack_7398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2950_delayed_1_0_3028_inst_ack_1, ack => convolve_CP_6745_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: 	156 
    -- CP-element group 214: 	188 
    -- CP-element group 214: 	172 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_Sample/req
      -- 
    req_7406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(214), ack => WPIPE_xxconvolvexxconv_ip4_3032_inst_req_0); -- 
    convolve_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(213) & convolve_CP_6745_elements(156) & convolve_CP_6745_elements(188) & convolve_CP_6745_elements(172) & convolve_CP_6745_elements(216);
      gj_convolve_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	154 
    -- CP-element group 215: 	186 
    -- CP-element group 215: 	211 
    -- CP-element group 215: 	170 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_update_start_
      -- CP-element group 215: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_Update/req
      -- 
    ack_7407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip4_3032_inst_ack_0, ack => convolve_CP_6745_elements(215)); -- 
    req_7411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(215), ack => WPIPE_xxconvolvexxconv_ip4_3032_inst_req_1); -- 
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	317 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_ip4_3032_Update/ack
      -- 
    ack_7412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip4_3032_inst_ack_1, ack => convolve_CP_6745_elements(216)); -- 
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	23 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	220 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_sample_start_
      -- CP-element group 217: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_Sample/$entry
      -- CP-element group 217: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_Sample/rr
      -- 
    rr_7420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(217), ack => RPIPE_kernel_pipe1_3062_inst_req_0); -- 
    convolve_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(220);
      gj_convolve_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	219 
    -- CP-element group 218: 	89 
    -- CP-element group 218: 	70 
    -- CP-element group 218: 	26 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	300 
    -- CP-element group 218: 	311 
    -- CP-element group 218: 	270 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	85 
    -- CP-element group 218: 	66 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_update_start_
      -- CP-element group 218: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_Update/cr
      -- 
    cr_7425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(218), ack => RPIPE_kernel_pipe1_3062_inst_req_1); -- 
    convolve_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(219) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(270);
      gj_convolve_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	218 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_Sample/ra
      -- 
    ra_7421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_3062_inst_ack_0, ack => convolve_CP_6745_elements(219)); -- 
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	298 
    -- CP-element group 220: 	309 
    -- CP-element group 220: 	269 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	29 
    -- CP-element group 220: 	217 
    -- CP-element group 220: 	46 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe1_3062_Update/ca
      -- 
    ca_7426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_3062_inst_ack_1, ack => convolve_CP_6745_elements(220)); -- 
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	23 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	224 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_sample_start_
      -- CP-element group 221: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_Sample/rr
      -- 
    rr_7434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(221), ack => RPIPE_kernel_pipe2_3066_inst_req_0); -- 
    convolve_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(224);
      gj_convolve_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	89 
    -- CP-element group 222: 	70 
    -- CP-element group 222: 	26 
    -- CP-element group 222: 	223 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	300 
    -- CP-element group 222: 	311 
    -- CP-element group 222: 	277 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	85 
    -- CP-element group 222: 	66 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_update_start_
      -- CP-element group 222: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_Update/$entry
      -- CP-element group 222: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_Update/cr
      -- 
    cr_7439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(222), ack => RPIPE_kernel_pipe2_3066_inst_req_1); -- 
    convolve_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(223) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(277);
      gj_convolve_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	222 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_Sample/ra
      -- 
    ra_7435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_3066_inst_ack_0, ack => convolve_CP_6745_elements(223)); -- 
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	298 
    -- CP-element group 224: 	309 
    -- CP-element group 224: 	276 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	29 
    -- CP-element group 224: 	221 
    -- CP-element group 224: 	46 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe2_3066_Update/ca
      -- 
    ca_7440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_3066_inst_ack_1, ack => convolve_CP_6745_elements(224)); -- 
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	23 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	228 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_Sample/rr
      -- 
    rr_7448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(225), ack => RPIPE_kernel_pipe3_3070_inst_req_0); -- 
    convolve_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(228);
      gj_convolve_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	89 
    -- CP-element group 226: 	70 
    -- CP-element group 226: 	26 
    -- CP-element group 226: 	227 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	284 
    -- CP-element group 226: 	300 
    -- CP-element group 226: 	311 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	85 
    -- CP-element group 226: 	66 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_update_start_
      -- CP-element group 226: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_Update/cr
      -- 
    cr_7453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(226), ack => RPIPE_kernel_pipe3_3070_inst_req_1); -- 
    convolve_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(227) & convolve_CP_6745_elements(284) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311);
      gj_convolve_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	226 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_Sample/ra
      -- 
    ra_7449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_3070_inst_ack_0, ack => convolve_CP_6745_elements(227)); -- 
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	283 
    -- CP-element group 228: 	298 
    -- CP-element group 228: 	309 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	29 
    -- CP-element group 228: 	46 
    -- CP-element group 228: 	225 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_kernel_pipe3_3070_Update/ca
      -- 
    ca_7454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_3070_inst_ack_1, ack => convolve_CP_6745_elements(228)); -- 
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	23 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	232 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_Sample/rr
      -- 
    rr_7462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(229), ack => RPIPE_xxconvolvexxconv_k1_3074_inst_req_0); -- 
    convolve_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(232);
      gj_convolve_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	89 
    -- CP-element group 230: 	70 
    -- CP-element group 230: 	26 
    -- CP-element group 230: 	231 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	300 
    -- CP-element group 230: 	311 
    -- CP-element group 230: 	270 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	85 
    -- CP-element group 230: 	66 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_update_start_
      -- CP-element group 230: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_Update/cr
      -- 
    cr_7467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(230), ack => RPIPE_xxconvolvexxconv_k1_3074_inst_req_1); -- 
    convolve_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(231) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(270);
      gj_convolve_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	230 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_Sample/ra
      -- 
    ra_7463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_3074_inst_ack_0, ack => convolve_CP_6745_elements(231)); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	298 
    -- CP-element group 232: 	309 
    -- CP-element group 232: 	269 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	29 
    -- CP-element group 232: 	46 
    -- CP-element group 232: 	229 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k1_3074_Update/ca
      -- 
    ca_7468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_3074_inst_ack_1, ack => convolve_CP_6745_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	23 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	236 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_Sample/rr
      -- 
    rr_7476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(233), ack => RPIPE_xxconvolvexxconv_k2_3078_inst_req_0); -- 
    convolve_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(236);
      gj_convolve_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	89 
    -- CP-element group 234: 	70 
    -- CP-element group 234: 	26 
    -- CP-element group 234: 	235 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	300 
    -- CP-element group 234: 	311 
    -- CP-element group 234: 	277 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	85 
    -- CP-element group 234: 	66 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_update_start_
      -- CP-element group 234: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_Update/cr
      -- 
    cr_7481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(234), ack => RPIPE_xxconvolvexxconv_k2_3078_inst_req_1); -- 
    convolve_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(235) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(277);
      gj_convolve_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	234 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_Sample/ra
      -- 
    ra_7477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_3078_inst_ack_0, ack => convolve_CP_6745_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	298 
    -- CP-element group 236: 	309 
    -- CP-element group 236: 	276 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	29 
    -- CP-element group 236: 	46 
    -- CP-element group 236: 	233 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k2_3078_Update/ca
      -- 
    ca_7482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_3078_inst_ack_1, ack => convolve_CP_6745_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	23 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	240 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_Sample/rr
      -- 
    rr_7490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(237), ack => RPIPE_xxconvolvexxconv_k3_3082_inst_req_0); -- 
    convolve_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(240);
      gj_convolve_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: 	89 
    -- CP-element group 238: 	70 
    -- CP-element group 238: 	26 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	284 
    -- CP-element group 238: 	300 
    -- CP-element group 238: 	311 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	85 
    -- CP-element group 238: 	66 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_update_start_
      -- CP-element group 238: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_Update/cr
      -- 
    cr_7495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(238), ack => RPIPE_xxconvolvexxconv_k3_3082_inst_req_1); -- 
    convolve_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(239) & convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(284) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311);
      gj_convolve_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	238 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_Sample/ra
      -- 
    ra_7491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_3082_inst_ack_0, ack => convolve_CP_6745_elements(239)); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	283 
    -- CP-element group 240: 	298 
    -- CP-element group 240: 	309 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	29 
    -- CP-element group 240: 	237 
    -- CP-element group 240: 	46 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/RPIPE_xxconvolvexxconv_k3_3082_Update/ca
      -- 
    ca_7496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_3082_inst_ack_1, ack => convolve_CP_6745_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	89 
    -- CP-element group 241: 	70 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_Sample/req
      -- CP-element group 241: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_sample_start_
      -- 
    req_7504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(241), ack => W_read_k_3004_delayed_1_0_3084_inst_req_0); -- 
    convolve_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(243);
      gj_convolve_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	26 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	300 
    -- CP-element group 242: 	311 
    -- CP-element group 242: 	244 
    -- CP-element group 242: 	270 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_Update/req
      -- CP-element group 242: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_update_start_
      -- 
    req_7509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(242), ack => W_read_k_3004_delayed_1_0_3084_inst_req_1); -- 
    convolve_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(244) & convolve_CP_6745_elements(270);
      gj_convolve_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: 	85 
    -- CP-element group 243: 	66 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_sample_completed_
      -- 
    ack_7505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_3004_delayed_1_0_3084_inst_ack_0, ack => convolve_CP_6745_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	298 
    -- CP-element group 244: 	309 
    -- CP-element group 244: 	269 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	29 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	46 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3086_update_completed_
      -- 
    ack_7510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_3004_delayed_1_0_3084_inst_ack_1, ack => convolve_CP_6745_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	89 
    -- CP-element group 245: 	70 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_Sample/req
      -- CP-element group 245: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_sample_start_
      -- 
    req_7518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(245), ack => W_read_k_3010_delayed_1_0_3093_inst_req_0); -- 
    convolve_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(247);
      gj_convolve_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	26 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	300 
    -- CP-element group 246: 	311 
    -- CP-element group 246: 	248 
    -- CP-element group 246: 	277 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_Update/req
      -- CP-element group 246: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_update_start_
      -- 
    req_7523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(246), ack => W_read_k_3010_delayed_1_0_3093_inst_req_1); -- 
    convolve_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(248) & convolve_CP_6745_elements(277);
      gj_convolve_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: 	85 
    -- CP-element group 247: 	66 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_sample_completed_
      -- 
    ack_7519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_3010_delayed_1_0_3093_inst_ack_0, ack => convolve_CP_6745_elements(247)); -- 
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	298 
    -- CP-element group 248: 	309 
    -- CP-element group 248: 	276 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	29 
    -- CP-element group 248: 	246 
    -- CP-element group 248: 	46 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3095_Update/ack
      -- 
    ack_7524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_3010_delayed_1_0_3093_inst_ack_1, ack => convolve_CP_6745_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	89 
    -- CP-element group 249: 	70 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_Sample/req
      -- CP-element group 249: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_sample_start_
      -- 
    req_7532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(249), ack => W_read_k_3016_delayed_1_0_3102_inst_req_0); -- 
    convolve_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(251);
      gj_convolve_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	26 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	284 
    -- CP-element group 250: 	300 
    -- CP-element group 250: 	311 
    -- CP-element group 250: 	252 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_Update/req
      -- CP-element group 250: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_update_start_
      -- 
    req_7537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(250), ack => W_read_k_3016_delayed_1_0_3102_inst_req_1); -- 
    convolve_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(284) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(252);
      gj_convolve_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: 	85 
    -- CP-element group 251: 	66 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_sample_completed_
      -- 
    ack_7533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_3016_delayed_1_0_3102_inst_ack_0, ack => convolve_CP_6745_elements(251)); -- 
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	283 
    -- CP-element group 252: 	298 
    -- CP-element group 252: 	309 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	29 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	46 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3104_update_completed_
      -- 
    ack_7538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_3016_delayed_1_0_3102_inst_ack_1, ack => convolve_CP_6745_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	32 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_Sample/req
      -- CP-element group 253: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_sample_start_
      -- 
    req_7546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(253), ack => W_acc1_3070_delayed_1_0_3159_inst_req_0); -- 
    convolve_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(32) & convolve_CP_6745_elements(255);
      gj_convolve_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	26 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	300 
    -- CP-element group 254: 	256 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_Update/req
      -- CP-element group 254: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_update_start_
      -- 
    req_7551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(254), ack => W_acc1_3070_delayed_1_0_3159_inst_req_1); -- 
    convolve_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(256);
      gj_convolve_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	30 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_sample_completed_
      -- 
    ack_7547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc1_3070_delayed_1_0_3159_inst_ack_0, ack => convolve_CP_6745_elements(255)); -- 
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	298 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	29 
    -- CP-element group 256: 	254 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3161_update_completed_
      -- 
    ack_7552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc1_3070_delayed_1_0_3159_inst_ack_1, ack => convolve_CP_6745_elements(256)); -- 
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	51 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_Sample/req
      -- CP-element group 257: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_Sample/$entry
      -- CP-element group 257: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_sample_start_
      -- 
    req_7560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(257), ack => W_acc2_3079_delayed_1_0_3171_inst_req_0); -- 
    convolve_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(51) & convolve_CP_6745_elements(259);
      gj_convolve_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	26 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	311 
    -- CP-element group 258: 	260 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_Update/req
      -- CP-element group 258: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_update_start_
      -- 
    req_7565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(258), ack => W_acc2_3079_delayed_1_0_3171_inst_req_1); -- 
    convolve_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(260);
      gj_convolve_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: 	47 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_sample_completed_
      -- 
    ack_7561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc2_3079_delayed_1_0_3171_inst_ack_0, ack => convolve_CP_6745_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	309 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	46 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3173_update_completed_
      -- 
    ack_7566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc2_3079_delayed_1_0_3171_inst_ack_1, ack => convolve_CP_6745_elements(260)); -- 
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	23 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_Sample/rr
      -- CP-element group 261: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_sample_start_
      -- 
    rr_7574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(261), ack => SUB_u16_u16_3208_inst_req_0); -- 
    convolve_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(23) & convolve_CP_6745_elements(263);
      gj_convolve_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	281 
    -- CP-element group 262: 	264 
    -- CP-element group 262: 	267 
    -- CP-element group 262: 	274 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_update_start_
      -- 
    cr_7579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(262), ack => SUB_u16_u16_3208_inst_req_1); -- 
    convolve_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(281) & convolve_CP_6745_elements(264) & convolve_CP_6745_elements(267) & convolve_CP_6745_elements(274);
      gj_convolve_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_Sample/ra
      -- 
    ra_7575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3208_inst_ack_0, ack => convolve_CP_6745_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	24 
    -- CP-element group 264: 	265 
    -- CP-element group 264: 	272 
    -- CP-element group 264: 	279 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_Update/ca
      -- CP-element group 264: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/SUB_u16_u16_3208_update_completed_
      -- 
    ca_7580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3208_inst_ack_1, ack => convolve_CP_6745_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	89 
    -- CP-element group 265: 	70 
    -- CP-element group 265: 	264 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_Sample/req
      -- CP-element group 265: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_sample_start_
      -- 
    req_7588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(265), ack => W_store_kernel_3127_delayed_1_0_3226_inst_req_0); -- 
    convolve_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(264) & convolve_CP_6745_elements(267);
      gj_convolve_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: 	270 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_Update/req
      -- CP-element group 266: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_update_start_
      -- 
    req_7593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(266), ack => W_store_kernel_3127_delayed_1_0_3226_inst_req_1); -- 
    convolve_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(268) & convolve_CP_6745_elements(270);
      gj_convolve_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	262 
    -- CP-element group 267: 	85 
    -- CP-element group 267: 	66 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_Sample/$exit
      -- 
    ack_7589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_3127_delayed_1_0_3226_inst_ack_0, ack => convolve_CP_6745_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3228_update_completed_
      -- 
    ack_7594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_3127_delayed_1_0_3226_inst_ack_1, ack => convolve_CP_6745_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	220 
    -- CP-element group 269: 	244 
    -- CP-element group 269: 	232 
    -- CP-element group 269: 	268 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_Sample/req
      -- 
    req_7602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(269), ack => WPIPE_xxconvolvexxconv_k1_3230_inst_req_0); -- 
    convolve_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(220) & convolve_CP_6745_elements(244) & convolve_CP_6745_elements(232) & convolve_CP_6745_elements(268) & convolve_CP_6745_elements(271);
      gj_convolve_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	218 
    -- CP-element group 270: 	242 
    -- CP-element group 270: 	230 
    -- CP-element group 270: 	266 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_update_start_
      -- CP-element group 270: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_Update/req
      -- CP-element group 270: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_Sample/ack
      -- 
    ack_7603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_3230_inst_ack_0, ack => convolve_CP_6745_elements(270)); -- 
    req_7607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(270), ack => WPIPE_xxconvolvexxconv_k1_3230_inst_req_1); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	317 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k1_3230_Update/ack
      -- 
    ack_7608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_3230_inst_ack_1, ack => convolve_CP_6745_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	89 
    -- CP-element group 272: 	70 
    -- CP-element group 272: 	264 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_sample_start_
      -- 
    req_7616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(272), ack => W_store_kernel_3131_delayed_1_0_3233_inst_req_0); -- 
    convolve_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(264) & convolve_CP_6745_elements(274);
      gj_convolve_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: 	277 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_Update/req
      -- CP-element group 273: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_update_start_
      -- CP-element group 273: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_Update/$entry
      -- 
    req_7621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(273), ack => W_store_kernel_3131_delayed_1_0_3233_inst_req_1); -- 
    convolve_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(275) & convolve_CP_6745_elements(277);
      gj_convolve_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	262 
    -- CP-element group 274: 	85 
    -- CP-element group 274: 	66 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_Sample/ack
      -- CP-element group 274: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_Sample/$exit
      -- 
    ack_7617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_3131_delayed_1_0_3233_inst_ack_0, ack => convolve_CP_6745_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3235_Update/ack
      -- 
    ack_7622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_3131_delayed_1_0_3233_inst_ack_1, ack => convolve_CP_6745_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	236 
    -- CP-element group 276: 	248 
    -- CP-element group 276: 	224 
    -- CP-element group 276: 	275 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_sample_start_
      -- 
    req_7630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(276), ack => WPIPE_xxconvolvexxconv_k2_3237_inst_req_0); -- 
    convolve_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(236) & convolve_CP_6745_elements(248) & convolve_CP_6745_elements(224) & convolve_CP_6745_elements(275) & convolve_CP_6745_elements(278);
      gj_convolve_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	222 
    -- CP-element group 277: 	246 
    -- CP-element group 277: 	234 
    -- CP-element group 277: 	273 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_Update/req
      -- CP-element group 277: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_update_start_
      -- CP-element group 277: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_sample_completed_
      -- 
    ack_7631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_3237_inst_ack_0, ack => convolve_CP_6745_elements(277)); -- 
    req_7635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(277), ack => WPIPE_xxconvolvexxconv_k2_3237_inst_req_1); -- 
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	317 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k2_3237_update_completed_
      -- 
    ack_7636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_3237_inst_ack_1, ack => convolve_CP_6745_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	89 
    -- CP-element group 279: 	70 
    -- CP-element group 279: 	264 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_Sample/req
      -- CP-element group 279: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_Sample/$entry
      -- 
    req_7644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(279), ack => W_store_kernel_3135_delayed_1_0_3240_inst_req_0); -- 
    convolve_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(89) & convolve_CP_6745_elements(70) & convolve_CP_6745_elements(264) & convolve_CP_6745_elements(281);
      gj_convolve_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	282 
    -- CP-element group 280: 	284 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_update_start_
      -- CP-element group 280: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_Update/$entry
      -- CP-element group 280: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_Update/req
      -- 
    req_7649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(280), ack => W_store_kernel_3135_delayed_1_0_3240_inst_req_1); -- 
    convolve_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(282) & convolve_CP_6745_elements(284);
      gj_convolve_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281: marked-successors 
    -- CP-element group 281: 	262 
    -- CP-element group 281: 	85 
    -- CP-element group 281: 	66 
    -- CP-element group 281: 	279 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_Sample/ack
      -- 
    ack_7645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_3135_delayed_1_0_3240_inst_ack_0, ack => convolve_CP_6745_elements(281)); -- 
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3242_Update/ack
      -- 
    ack_7650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_3135_delayed_1_0_3240_inst_ack_1, ack => convolve_CP_6745_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: 	240 
    -- CP-element group 283: 	252 
    -- CP-element group 283: 	228 
    -- CP-element group 283: marked-predecessors 
    -- CP-element group 283: 	285 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_Sample/req
      -- 
    req_7658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(283), ack => WPIPE_xxconvolvexxconv_k3_3244_inst_req_0); -- 
    convolve_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(282) & convolve_CP_6745_elements(240) & convolve_CP_6745_elements(252) & convolve_CP_6745_elements(228) & convolve_CP_6745_elements(285);
      gj_convolve_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	238 
    -- CP-element group 284: 	250 
    -- CP-element group 284: 	226 
    -- CP-element group 284: 	280 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_update_start_
      -- CP-element group 284: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_Update/req
      -- 
    ack_7659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_3244_inst_ack_0, ack => convolve_CP_6745_elements(284)); -- 
    req_7663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(284), ack => WPIPE_xxconvolvexxconv_k3_3244_inst_req_1); -- 
    -- CP-element group 285:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	317 
    -- CP-element group 285: marked-successors 
    -- CP-element group 285: 	283 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_xxconvolvexxconv_k3_3244_Update/ack
      -- 
    ack_7664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_3244_inst_ack_1, ack => convolve_CP_6745_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	108 
    -- CP-element group 286: 	127 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	288 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_Sample/req
      -- 
    req_7672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(286), ack => W_num_done_3178_delayed_1_0_3285_inst_req_0); -- 
    convolve_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(127) & convolve_CP_6745_elements(288);
      gj_convolve_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	26 
    -- CP-element group 287: marked-predecessors 
    -- CP-element group 287: 	289 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	289 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_update_start_
      -- CP-element group 287: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_Update/req
      -- 
    req_7677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(287), ack => W_num_done_3178_delayed_1_0_3285_inst_req_1); -- 
    convolve_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(289);
      gj_convolve_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: 	104 
    -- CP-element group 288: 	123 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_Sample/ack
      -- 
    ack_7673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3178_delayed_1_0_3285_inst_ack_0, ack => convolve_CP_6745_elements(288)); -- 
    -- CP-element group 289:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	317 
    -- CP-element group 289: marked-successors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: 	29 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3287_Update/ack
      -- 
    ack_7678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3178_delayed_1_0_3285_inst_ack_1, ack => convolve_CP_6745_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	108 
    -- CP-element group 290: 	127 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_Sample/req
      -- 
    req_7686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(290), ack => W_num_done_3184_delayed_1_0_3294_inst_req_0); -- 
    convolve_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(127) & convolve_CP_6745_elements(292);
      gj_convolve_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	26 
    -- CP-element group 291: marked-predecessors 
    -- CP-element group 291: 	293 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_update_start_
      -- CP-element group 291: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_Update/req
      -- 
    req_7691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(291), ack => W_num_done_3184_delayed_1_0_3294_inst_req_1); -- 
    convolve_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(26) & convolve_CP_6745_elements(293);
      gj_convolve_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: 	104 
    -- CP-element group 292: 	123 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_Sample/ack
      -- 
    ack_7687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3184_delayed_1_0_3294_inst_ack_0, ack => convolve_CP_6745_elements(292)); -- 
    -- CP-element group 293:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	317 
    -- CP-element group 293: marked-successors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: 	46 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3296_Update/ack
      -- 
    ack_7692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3184_delayed_1_0_3294_inst_ack_1, ack => convolve_CP_6745_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	108 
    -- CP-element group 294: 	127 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_Sample/req
      -- 
    req_7700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(294), ack => W_num_done_3189_delayed_1_0_3303_inst_req_0); -- 
    convolve_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(127) & convolve_CP_6745_elements(296);
      gj_convolve_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: marked-predecessors 
    -- CP-element group 295: 	297 
    -- CP-element group 295: 	300 
    -- CP-element group 295: 	303 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	297 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_update_start_
      -- CP-element group 295: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_Update/req
      -- 
    req_7705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(295), ack => W_num_done_3189_delayed_1_0_3303_inst_req_1); -- 
    convolve_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(297) & convolve_CP_6745_elements(300) & convolve_CP_6745_elements(303);
      gj_convolve_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: 	104 
    -- CP-element group 296: 	123 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_sample_completed_
      -- CP-element group 296: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_Sample/ack
      -- 
    ack_7701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3189_delayed_1_0_3303_inst_ack_0, ack => convolve_CP_6745_elements(296)); -- 
    -- CP-element group 297:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	295 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297: 	302 
    -- CP-element group 297: marked-successors 
    -- CP-element group 297: 	295 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_update_completed_
      -- CP-element group 297: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3305_Update/ack
      -- 
    ack_7706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3189_delayed_1_0_3303_inst_ack_1, ack => convolve_CP_6745_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	164 
    -- CP-element group 298: 	148 
    -- CP-element group 298: 	152 
    -- CP-element group 298: 	297 
    -- CP-element group 298: 	220 
    -- CP-element group 298: 	144 
    -- CP-element group 298: 	236 
    -- CP-element group 298: 	240 
    -- CP-element group 298: 	244 
    -- CP-element group 298: 	248 
    -- CP-element group 298: 	252 
    -- CP-element group 298: 	256 
    -- CP-element group 298: 	180 
    -- CP-element group 298: 	184 
    -- CP-element group 298: 	176 
    -- CP-element group 298: 	160 
    -- CP-element group 298: 	168 
    -- CP-element group 298: 	224 
    -- CP-element group 298: 	228 
    -- CP-element group 298: 	232 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_Sample/rr
      -- 
    rr_7714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(298), ack => type_cast_3309_inst_req_0); -- 
    convolve_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(164) & convolve_CP_6745_elements(148) & convolve_CP_6745_elements(152) & convolve_CP_6745_elements(297) & convolve_CP_6745_elements(220) & convolve_CP_6745_elements(144) & convolve_CP_6745_elements(236) & convolve_CP_6745_elements(240) & convolve_CP_6745_elements(244) & convolve_CP_6745_elements(248) & convolve_CP_6745_elements(252) & convolve_CP_6745_elements(256) & convolve_CP_6745_elements(180) & convolve_CP_6745_elements(184) & convolve_CP_6745_elements(176) & convolve_CP_6745_elements(160) & convolve_CP_6745_elements(168) & convolve_CP_6745_elements(224) & convolve_CP_6745_elements(228) & convolve_CP_6745_elements(232) & convolve_CP_6745_elements(300);
      gj_convolve_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: marked-predecessors 
    -- CP-element group 299: 	301 
    -- CP-element group 299: 	303 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	301 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_update_start_
      -- CP-element group 299: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_Update/cr
      -- 
    cr_7719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(299), ack => type_cast_3309_inst_req_1); -- 
    convolve_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(301) & convolve_CP_6745_elements(303);
      gj_convolve_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	162 
    -- CP-element group 300: 	166 
    -- CP-element group 300: 	150 
    -- CP-element group 300: 	295 
    -- CP-element group 300: 	298 
    -- CP-element group 300: 	218 
    -- CP-element group 300: 	222 
    -- CP-element group 300: 	146 
    -- CP-element group 300: 	238 
    -- CP-element group 300: 	242 
    -- CP-element group 300: 	246 
    -- CP-element group 300: 	250 
    -- CP-element group 300: 	254 
    -- CP-element group 300: 	182 
    -- CP-element group 300: 	174 
    -- CP-element group 300: 	178 
    -- CP-element group 300: 	158 
    -- CP-element group 300: 	142 
    -- CP-element group 300: 	226 
    -- CP-element group 300: 	230 
    -- CP-element group 300: 	234 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_Sample/ra
      -- 
    ra_7715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3309_inst_ack_0, ack => convolve_CP_6745_elements(300)); -- 
    -- CP-element group 301:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	299 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301: marked-successors 
    -- CP-element group 301: 	299 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3309_Update/ca
      -- 
    ca_7720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3309_inst_ack_1, ack => convolve_CP_6745_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	297 
    -- CP-element group 302: 	301 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: 	315 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_Sample/req
      -- 
    req_7728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(302), ack => WPIPE_output_pipe_3307_inst_req_0); -- 
    convolve_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(297) & convolve_CP_6745_elements(301) & convolve_CP_6745_elements(304) & convolve_CP_6745_elements(315);
      gj_convolve_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	295 
    -- CP-element group 303: 	299 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_update_start_
      -- CP-element group 303: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_Update/req
      -- 
    ack_7729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3307_inst_ack_0, ack => convolve_CP_6745_elements(303)); -- 
    req_7733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(303), ack => WPIPE_output_pipe_3307_inst_req_1); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	313 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3307_Update/ack
      -- 
    ack_7734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3307_inst_ack_1, ack => convolve_CP_6745_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	108 
    -- CP-element group 305: 	127 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_Sample/req
      -- 
    req_7742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(305), ack => W_num_done_3194_delayed_1_0_3311_inst_req_0); -- 
    convolve_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(108) & convolve_CP_6745_elements(127) & convolve_CP_6745_elements(307);
      gj_convolve_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: 	311 
    -- CP-element group 306: 	314 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_update_start_
      -- CP-element group 306: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_Update/req
      -- 
    req_7747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(306), ack => W_num_done_3194_delayed_1_0_3311_inst_req_1); -- 
    convolve_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(308) & convolve_CP_6745_elements(311) & convolve_CP_6745_elements(314);
      gj_convolve_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	104 
    -- CP-element group 307: 	123 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_Sample/ack
      -- 
    ack_7743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3194_delayed_1_0_3311_inst_ack_0, ack => convolve_CP_6745_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308: 	313 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/assign_stmt_3313_Update/ack
      -- 
    ack_7748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3194_delayed_1_0_3311_inst_ack_1, ack => convolve_CP_6745_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	164 
    -- CP-element group 309: 	148 
    -- CP-element group 309: 	152 
    -- CP-element group 309: 	308 
    -- CP-element group 309: 	220 
    -- CP-element group 309: 	236 
    -- CP-element group 309: 	240 
    -- CP-element group 309: 	244 
    -- CP-element group 309: 	248 
    -- CP-element group 309: 	252 
    -- CP-element group 309: 	260 
    -- CP-element group 309: 	180 
    -- CP-element group 309: 	184 
    -- CP-element group 309: 	156 
    -- CP-element group 309: 	188 
    -- CP-element group 309: 	168 
    -- CP-element group 309: 	172 
    -- CP-element group 309: 	224 
    -- CP-element group 309: 	228 
    -- CP-element group 309: 	232 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_Sample/rr
      -- 
    rr_7756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(309), ack => type_cast_3317_inst_req_0); -- 
    convolve_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(164) & convolve_CP_6745_elements(148) & convolve_CP_6745_elements(152) & convolve_CP_6745_elements(308) & convolve_CP_6745_elements(220) & convolve_CP_6745_elements(236) & convolve_CP_6745_elements(240) & convolve_CP_6745_elements(244) & convolve_CP_6745_elements(248) & convolve_CP_6745_elements(252) & convolve_CP_6745_elements(260) & convolve_CP_6745_elements(180) & convolve_CP_6745_elements(184) & convolve_CP_6745_elements(156) & convolve_CP_6745_elements(188) & convolve_CP_6745_elements(168) & convolve_CP_6745_elements(172) & convolve_CP_6745_elements(224) & convolve_CP_6745_elements(228) & convolve_CP_6745_elements(232) & convolve_CP_6745_elements(311);
      gj_convolve_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	314 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_update_start_
      -- CP-element group 310: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_Update/cr
      -- 
    cr_7761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(310), ack => type_cast_3317_inst_req_1); -- 
    convolve_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(312) & convolve_CP_6745_elements(314);
      gj_convolve_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	162 
    -- CP-element group 311: 	166 
    -- CP-element group 311: 	150 
    -- CP-element group 311: 	154 
    -- CP-element group 311: 	306 
    -- CP-element group 311: 	309 
    -- CP-element group 311: 	218 
    -- CP-element group 311: 	222 
    -- CP-element group 311: 	146 
    -- CP-element group 311: 	238 
    -- CP-element group 311: 	242 
    -- CP-element group 311: 	246 
    -- CP-element group 311: 	250 
    -- CP-element group 311: 	258 
    -- CP-element group 311: 	182 
    -- CP-element group 311: 	186 
    -- CP-element group 311: 	178 
    -- CP-element group 311: 	170 
    -- CP-element group 311: 	226 
    -- CP-element group 311: 	230 
    -- CP-element group 311: 	234 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_Sample/ra
      -- 
    ra_7757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3317_inst_ack_0, ack => convolve_CP_6745_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/type_cast_3317_Update/ca
      -- 
    ca_7762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3317_inst_ack_1, ack => convolve_CP_6745_elements(312)); -- 
    -- CP-element group 313:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	304 
    -- CP-element group 313: 	308 
    -- CP-element group 313: 	312 
    -- CP-element group 313: marked-predecessors 
    -- CP-element group 313: 	315 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_Sample/req
      -- 
    req_7770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(313), ack => WPIPE_output_pipe_3315_inst_req_0); -- 
    convolve_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(304) & convolve_CP_6745_elements(308) & convolve_CP_6745_elements(312) & convolve_CP_6745_elements(315);
      gj_convolve_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	306 
    -- CP-element group 314: 	310 
    -- CP-element group 314:  members (6) 
      -- CP-element group 314: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_sample_completed_
      -- CP-element group 314: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_update_start_
      -- CP-element group 314: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_Sample/ack
      -- CP-element group 314: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_Update/$entry
      -- CP-element group 314: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_Update/req
      -- 
    ack_7771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3315_inst_ack_0, ack => convolve_CP_6745_elements(314)); -- 
    req_7775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(314), ack => WPIPE_output_pipe_3315_inst_req_1); -- 
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	302 
    -- CP-element group 315: 	313 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_update_completed_
      -- CP-element group 315: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_Update/$exit
      -- CP-element group 315: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/WPIPE_output_pipe_3315_Update/ack
      -- 
    ack_7776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3315_inst_ack_1, ack => convolve_CP_6745_elements(315)); -- 
    -- CP-element group 316:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	23 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	24 
    -- CP-element group 316:  members (1) 
      -- CP-element group 316: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_6745_elements(316) is a control-delay.
    cp_element_316_delay: control_delay_element  generic map(name => " 316_delay", delay_value => 1)  port map(req => convolve_CP_6745_elements(23), ack => convolve_CP_6745_elements(316), clk => clk, reset =>reset);
    -- CP-element group 317:  join  transition  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	285 
    -- CP-element group 317: 	289 
    -- CP-element group 317: 	293 
    -- CP-element group 317: 	315 
    -- CP-element group 317: 	216 
    -- CP-element group 317: 	202 
    -- CP-element group 317: 	26 
    -- CP-element group 317: 	209 
    -- CP-element group 317: 	195 
    -- CP-element group 317: 	271 
    -- CP-element group 317: 	278 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	20 
    -- CP-element group 317:  members (1) 
      -- CP-element group 317: 	 branch_block_stmt_2870/do_while_stmt_2887/do_while_stmt_2887_loop_body/$exit
      -- 
    convolve_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolve_CP_6745_elements(285) & convolve_CP_6745_elements(289) & convolve_CP_6745_elements(293) & convolve_CP_6745_elements(315) & convolve_CP_6745_elements(216) & convolve_CP_6745_elements(202) & convolve_CP_6745_elements(26) & convolve_CP_6745_elements(209) & convolve_CP_6745_elements(195) & convolve_CP_6745_elements(271) & convolve_CP_6745_elements(278);
      gj_convolve_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6745_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	19 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_2870/do_while_stmt_2887/loop_exit/$exit
      -- CP-element group 318: 	 branch_block_stmt_2870/do_while_stmt_2887/loop_exit/ack
      -- 
    ack_7781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2887_branch_ack_0, ack => convolve_CP_6745_elements(318)); -- 
    -- CP-element group 319:  transition  input  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	19 
    -- CP-element group 319: successors 
    -- CP-element group 319:  members (2) 
      -- CP-element group 319: 	 branch_block_stmt_2870/do_while_stmt_2887/loop_taken/$exit
      -- CP-element group 319: 	 branch_block_stmt_2870/do_while_stmt_2887/loop_taken/ack
      -- 
    ack_7785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2887_branch_ack_1, ack => convolve_CP_6745_elements(319)); -- 
    -- CP-element group 320:  transition  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	17 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	2 
    -- CP-element group 320:  members (1) 
      -- CP-element group 320: 	 branch_block_stmt_2870/do_while_stmt_2887/$exit
      -- 
    convolve_CP_6745_elements(320) <= convolve_CP_6745_elements(17);
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	2 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_sample_completed_
      -- CP-element group 321: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_update_start_
      -- CP-element group 321: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_Sample/ack
      -- CP-element group 321: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_Update/req
      -- 
    ack_7798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3322_inst_ack_0, ack => convolve_CP_6745_elements(321)); -- 
    req_7802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(321), ack => WPIPE_input_done_pipe_3322_inst_req_1); -- 
    -- CP-element group 322:  transition  place  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (8) 
      -- CP-element group 322: 	 branch_block_stmt_2870/loopback
      -- CP-element group 322: 	 branch_block_stmt_2870/assign_stmt_3324__exit__
      -- CP-element group 322: 	 branch_block_stmt_2870/assign_stmt_3324/$exit
      -- CP-element group 322: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_update_completed_
      -- CP-element group 322: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_2870/assign_stmt_3324/WPIPE_input_done_pipe_3322_Update/ack
      -- CP-element group 322: 	 branch_block_stmt_2870/loopback_PhiReq/$entry
      -- CP-element group 322: 	 branch_block_stmt_2870/loopback_PhiReq/$exit
      -- 
    ack_7803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3322_inst_ack_1, ack => convolve_CP_6745_elements(322)); -- 
    -- CP-element group 323:  merge  fork  transition  place  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	0 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	6 
    -- CP-element group 323: 	10 
    -- CP-element group 323: 	11 
    -- CP-element group 323: 	14 
    -- CP-element group 323: 	3 
    -- CP-element group 323:  members (22) 
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_update_start_
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_Sample/rr
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_size_pipe_2883_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_Update/cr
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_Sample/rr
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_update_start_
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2880_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_Update/cr
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/RPIPE_num_out_pipe_2873_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_Update/cr
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886__entry__
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2875_update_start_
      -- CP-element group 323: 	 branch_block_stmt_2870/merge_stmt_2871__exit__
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/$entry
      -- CP-element group 323: 	 branch_block_stmt_2870/assign_stmt_2876_to_assign_stmt_2886/SUB_u16_u16_2885_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_2870/merge_stmt_2871_PhiReqMerge
      -- CP-element group 323: 	 branch_block_stmt_2870/merge_stmt_2871_PhiAck/$entry
      -- CP-element group 323: 	 branch_block_stmt_2870/merge_stmt_2871_PhiAck/$exit
      -- CP-element group 323: 	 branch_block_stmt_2870/merge_stmt_2871_PhiAck/dummy
      -- 
    rr_6832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(323), ack => RPIPE_size_pipe_2883_inst_req_0); -- 
    cr_6819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(323), ack => SUB_u16_u16_2880_inst_req_1); -- 
    rr_6776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(323), ack => RPIPE_num_out_pipe_2873_inst_req_0); -- 
    cr_6791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(323), ack => SUB_u16_u16_2875_inst_req_1); -- 
    cr_6847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6745_elements(323), ack => SUB_u16_u16_2885_inst_req_1); -- 
    convolve_CP_6745_elements(323) <= OrReduce(convolve_CP_6745_elements(0) & convolve_CP_6745_elements(322));
    convolve_do_while_stmt_2887_terminator_7786: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_2887_terminator_7786", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_6745_elements(20),loop_continue => convolve_CP_6745_elements(319),loop_terminate => convolve_CP_6745_elements(318),loop_back => convolve_CP_6745_elements(18),loop_exit => convolve_CP_6745_elements(17),clk => clk, reset => reset); -- 
    phi_stmt_2889_phi_seq_6912_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6745_elements(35);
      convolve_CP_6745_elements(38)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6745_elements(38);
      convolve_CP_6745_elements(39)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6745_elements(40);
      convolve_CP_6745_elements(36) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6745_elements(33);
      convolve_CP_6745_elements(42)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6745_elements(44);
      convolve_CP_6745_elements(43)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6745_elements(45);
      convolve_CP_6745_elements(34) <= phi_mux_reqs(1);
      phi_stmt_2889_phi_seq_6912 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2889_phi_seq_6912") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6745_elements(25), 
          phi_sample_ack => convolve_CP_6745_elements(31), 
          phi_update_req => convolve_CP_6745_elements(27), 
          phi_update_ack => convolve_CP_6745_elements(32), 
          phi_mux_ack => convolve_CP_6745_elements(37), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2895_phi_seq_6956_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6745_elements(54);
      convolve_CP_6745_elements(57)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6745_elements(57);
      convolve_CP_6745_elements(58)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6745_elements(59);
      convolve_CP_6745_elements(55) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6745_elements(52);
      convolve_CP_6745_elements(61)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6745_elements(63);
      convolve_CP_6745_elements(62)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6745_elements(64);
      convolve_CP_6745_elements(53) <= phi_mux_reqs(1);
      phi_stmt_2895_phi_seq_6956 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2895_phi_seq_6956") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6745_elements(48), 
          phi_sample_ack => convolve_CP_6745_elements(49), 
          phi_update_req => convolve_CP_6745_elements(50), 
          phi_update_ack => convolve_CP_6745_elements(51), 
          phi_mux_ack => convolve_CP_6745_elements(56), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2900_phi_seq_7000_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6745_elements(73);
      convolve_CP_6745_elements(76)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6745_elements(76);
      convolve_CP_6745_elements(77)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6745_elements(78);
      convolve_CP_6745_elements(74) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6745_elements(71);
      convolve_CP_6745_elements(80)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6745_elements(82);
      convolve_CP_6745_elements(81)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6745_elements(83);
      convolve_CP_6745_elements(72) <= phi_mux_reqs(1);
      phi_stmt_2900_phi_seq_7000 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2900_phi_seq_7000") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6745_elements(67), 
          phi_sample_ack => convolve_CP_6745_elements(68), 
          phi_update_req => convolve_CP_6745_elements(69), 
          phi_update_ack => convolve_CP_6745_elements(70), 
          phi_mux_ack => convolve_CP_6745_elements(75), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2905_phi_seq_7044_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6745_elements(92);
      convolve_CP_6745_elements(95)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6745_elements(95);
      convolve_CP_6745_elements(96)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6745_elements(97);
      convolve_CP_6745_elements(93) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6745_elements(90);
      convolve_CP_6745_elements(99)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6745_elements(101);
      convolve_CP_6745_elements(100)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6745_elements(102);
      convolve_CP_6745_elements(91) <= phi_mux_reqs(1);
      phi_stmt_2905_phi_seq_7044 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2905_phi_seq_7044") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6745_elements(86), 
          phi_sample_ack => convolve_CP_6745_elements(87), 
          phi_update_req => convolve_CP_6745_elements(88), 
          phi_update_ack => convolve_CP_6745_elements(89), 
          phi_mux_ack => convolve_CP_6745_elements(94), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2910_phi_seq_7088_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6745_elements(111);
      convolve_CP_6745_elements(114)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6745_elements(114);
      convolve_CP_6745_elements(115)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6745_elements(116);
      convolve_CP_6745_elements(112) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6745_elements(109);
      convolve_CP_6745_elements(118)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6745_elements(120);
      convolve_CP_6745_elements(119)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6745_elements(121);
      convolve_CP_6745_elements(110) <= phi_mux_reqs(1);
      phi_stmt_2910_phi_seq_7088 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2910_phi_seq_7088") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6745_elements(105), 
          phi_sample_ack => convolve_CP_6745_elements(106), 
          phi_update_req => convolve_CP_6745_elements(107), 
          phi_update_ack => convolve_CP_6745_elements(108), 
          phi_mux_ack => convolve_CP_6745_elements(113), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2915_phi_seq_7132_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6745_elements(130);
      convolve_CP_6745_elements(133)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6745_elements(133);
      convolve_CP_6745_elements(134)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6745_elements(135);
      convolve_CP_6745_elements(131) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6745_elements(128);
      convolve_CP_6745_elements(137)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6745_elements(139);
      convolve_CP_6745_elements(138)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6745_elements(140);
      convolve_CP_6745_elements(129) <= phi_mux_reqs(1);
      phi_stmt_2915_phi_seq_7132 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2915_phi_seq_7132") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6745_elements(124), 
          phi_sample_ack => convolve_CP_6745_elements(125), 
          phi_update_req => convolve_CP_6745_elements(126), 
          phi_update_ack => convolve_CP_6745_elements(127), 
          phi_mux_ack => convolve_CP_6745_elements(132), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6864_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_6745_elements(21);
        preds(1)  <= convolve_CP_6745_elements(22);
        entry_tmerge_6864 : transition_merge -- 
          generic map(name => " entry_tmerge_6864")
          port map (preds => preds, symbol_out => convolve_CP_6745_elements(23));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_i16_i16_3165_wire : std_logic_vector(15 downto 0);
    signal ADD_i16_i16_3168_wire : std_logic_vector(15 downto 0);
    signal ADD_i16_i16_3177_wire : std_logic_vector(15 downto 0);
    signal ADD_i16_i16_3180_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3252_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3272_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3281_wire : std_logic_vector(15 downto 0);
    signal ADD_u2_u2_3261_wire : std_logic_vector(1 downto 0);
    signal AND_u1_u1_3218_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2924_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_3054_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_3057_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2927_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3191_wire : std_logic_vector(0 downto 0);
    signal MUL_i16_i16_3126_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_3132_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_3138_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_3144_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_3150_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_3156_wire : std_logic_vector(15 downto 0);
    signal MUX_3262_wire : std_logic_vector(1 downto 0);
    signal MUX_3273_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_3321_wire : std_logic_vector(0 downto 0);
    signal RPIPE_num_out_pipe_2873_wire : std_logic_vector(15 downto 0);
    signal RPIPE_num_out_pipe_2878_wire : std_logic_vector(15 downto 0);
    signal RPIPE_size_pipe_2883_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_3113_3113_delayed_1_0_3209 : std_logic_vector(15 downto 0);
    signal UGT_u2_u1_3004_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_3001_wire : std_logic_vector(0 downto 0);
    signal acc1_2889 : std_logic_vector(15 downto 0);
    signal acc1_3070_delayed_1_0_3161 : std_logic_vector(15 downto 0);
    signal acc2_2895 : std_logic_vector(15 downto 0);
    signal acc2_3079_delayed_1_0_3173 : std_logic_vector(15 downto 0);
    signal acc_val1_3170 : std_logic_vector(15 downto 0);
    signal acc_val2_3182 : std_logic_vector(15 downto 0);
    signal all_done_flag_3225 : std_logic_vector(0 downto 0);
    signal chl_2915 : std_logic_vector(15 downto 0);
    signal chl_done_3187 : std_logic_vector(0 downto 0);
    signal col_2905 : std_logic_vector(15 downto 0);
    signal col_done_3199 : std_logic_vector(0 downto 0);
    signal iread1_2970 : std_logic_vector(15 downto 0);
    signal iread2_2979 : std_logic_vector(15 downto 0);
    signal iread3_2988 : std_logic_vector(15 downto 0);
    signal iread4_2997 : std_logic_vector(15 downto 0);
    signal ival1_3038 : std_logic_vector(15 downto 0);
    signal ival2_3042 : std_logic_vector(15 downto 0);
    signal ival3_3046 : std_logic_vector(15 downto 0);
    signal ival4_3050 : std_logic_vector(15 downto 0);
    signal konst_2874_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2879_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2884_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2923_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2926_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3003_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3053_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3056_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3190_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3207_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3249_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3251_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3258_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3260_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3269_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3271_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3280_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3290_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3299_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3323_wire_constant : std_logic_vector(7 downto 0);
    signal kread1_3092 : std_logic_vector(15 downto 0);
    signal kread2_3101 : std_logic_vector(15 downto 0);
    signal kread3_3110 : std_logic_vector(15 downto 0);
    signal kval1_3114 : std_logic_vector(15 downto 0);
    signal kval2_3118 : std_logic_vector(15 downto 0);
    signal kval3_3122 : std_logic_vector(15 downto 0);
    signal mul_val1_3128 : std_logic_vector(15 downto 0);
    signal mul_val2_3134 : std_logic_vector(15 downto 0);
    signal mul_val3_3140 : std_logic_vector(15 downto 0);
    signal mul_val4_3146 : std_logic_vector(15 downto 0);
    signal mul_val5_3152 : std_logic_vector(15 downto 0);
    signal mul_val6_3158 : std_logic_vector(15 downto 0);
    signal n_chl_3254 : std_logic_vector(15 downto 0);
    signal n_chl_3254_2919_buffered : std_logic_vector(15 downto 0);
    signal n_col_3276 : std_logic_vector(15 downto 0);
    signal n_col_3276_2909_buffered : std_logic_vector(15 downto 0);
    signal n_num_3265 : std_logic_vector(1 downto 0);
    signal n_num_3265_2914_buffered : std_logic_vector(1 downto 0);
    signal n_row_3284 : std_logic_vector(15 downto 0);
    signal n_row_3284_2904_buffered : std_logic_vector(15 downto 0);
    signal nacc1_3293 : std_logic_vector(15 downto 0);
    signal nacc1_3293_2894_buffered : std_logic_vector(15 downto 0);
    signal nacc2_3302 : std_logic_vector(15 downto 0);
    signal nacc2_3302_2899_buffered : std_logic_vector(15 downto 0);
    signal num_2910 : std_logic_vector(1 downto 0);
    signal num_chl_2886 : std_logic_vector(15 downto 0);
    signal num_col_2881 : std_logic_vector(15 downto 0);
    signal num_done_3178_delayed_1_0_3287 : std_logic_vector(0 downto 0);
    signal num_done_3184_delayed_1_0_3296 : std_logic_vector(0 downto 0);
    signal num_done_3189_delayed_1_0_3305 : std_logic_vector(0 downto 0);
    signal num_done_3194 : std_logic_vector(0 downto 0);
    signal num_done_3194_delayed_1_0_3313 : std_logic_vector(0 downto 0);
    signal num_row_2876 : std_logic_vector(15 downto 0);
    signal out_done_flag_3214 : std_logic_vector(0 downto 0);
    signal read_ip_2906_delayed_1_0_2964 : std_logic_vector(0 downto 0);
    signal read_ip_2912_delayed_1_0_2973 : std_logic_vector(0 downto 0);
    signal read_ip_2918_delayed_1_0_2982 : std_logic_vector(0 downto 0);
    signal read_ip_2924_delayed_1_0_2991 : std_logic_vector(0 downto 0);
    signal read_ip_2929 : std_logic_vector(0 downto 0);
    signal read_k_3004_delayed_1_0_3086 : std_logic_vector(0 downto 0);
    signal read_k_3010_delayed_1_0_3095 : std_logic_vector(0 downto 0);
    signal read_k_3016_delayed_1_0_3104 : std_logic_vector(0 downto 0);
    signal read_k_3059 : std_logic_vector(0 downto 0);
    signal row_2900 : std_logic_vector(15 downto 0);
    signal row_done_3204 : std_logic_vector(0 downto 0);
    signal store_kernel_3127_delayed_1_0_3228 : std_logic_vector(0 downto 0);
    signal store_kernel_3131_delayed_1_0_3235 : std_logic_vector(0 downto 0);
    signal store_kernel_3135_delayed_1_0_3242 : std_logic_vector(0 downto 0);
    signal store_kernel_3220 : std_logic_vector(0 downto 0);
    signal temp1_1_2949 : std_logic_vector(15 downto 0);
    signal temp1_2_2953 : std_logic_vector(15 downto 0);
    signal temp1_3_2957 : std_logic_vector(15 downto 0);
    signal temp1_4_2961 : std_logic_vector(15 downto 0);
    signal temp2_1_2933 : std_logic_vector(15 downto 0);
    signal temp2_2_2937 : std_logic_vector(15 downto 0);
    signal temp2_3_2941 : std_logic_vector(15 downto 0);
    signal temp2_4_2945 : std_logic_vector(15 downto 0);
    signal tempk1_1_3063 : std_logic_vector(15 downto 0);
    signal tempk1_2_3067 : std_logic_vector(15 downto 0);
    signal tempk1_3_3071 : std_logic_vector(15 downto 0);
    signal tempk2_1_3075 : std_logic_vector(15 downto 0);
    signal tempk2_2_3079 : std_logic_vector(15 downto 0);
    signal tempk2_3_3083 : std_logic_vector(15 downto 0);
    signal type_cast_2893_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2898_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2903_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2908_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2913_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_2918_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3309_wire : std_logic_vector(15 downto 0);
    signal type_cast_3317_wire : std_logic_vector(15 downto 0);
    signal write_input_2938_delayed_1_0_3009 : std_logic_vector(0 downto 0);
    signal write_input_2942_delayed_1_0_3016 : std_logic_vector(0 downto 0);
    signal write_input_2946_delayed_1_0_3023 : std_logic_vector(0 downto 0);
    signal write_input_2950_delayed_1_0_3030 : std_logic_vector(0 downto 0);
    signal write_input_3006 : std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip4
    signal xxconvolvexxconv_ip4_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip4_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip4_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip4
    signal xxconvolvexxconv_ip4_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip4_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip4_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_2874_wire_constant <= "0000000000000001";
    konst_2879_wire_constant <= "0000000000000001";
    konst_2884_wire_constant <= "0000000000000001";
    konst_2923_wire_constant <= "0000000000000000";
    konst_2926_wire_constant <= "10";
    konst_3003_wire_constant <= "00";
    konst_3053_wire_constant <= "0000000000000000";
    konst_3056_wire_constant <= "0000000000000000";
    konst_3190_wire_constant <= "10";
    konst_3207_wire_constant <= "0000000000000001";
    konst_3249_wire_constant <= "0000000000000000";
    konst_3251_wire_constant <= "0000000000000001";
    konst_3258_wire_constant <= "00";
    konst_3260_wire_constant <= "01";
    konst_3269_wire_constant <= "0000000000000000";
    konst_3271_wire_constant <= "0000000000000001";
    konst_3280_wire_constant <= "0000000000000010";
    konst_3290_wire_constant <= "0000000000000000";
    konst_3299_wire_constant <= "0000000000000000";
    konst_3323_wire_constant <= "00000001";
    type_cast_2893_wire_constant <= "0000000000000000";
    type_cast_2898_wire_constant <= "0000000000000000";
    type_cast_2903_wire_constant <= "0000000000000000";
    type_cast_2908_wire_constant <= "0000000000000000";
    type_cast_2913_wire_constant <= "00";
    type_cast_2918_wire_constant <= "0000000000000000";
    phi_stmt_2889: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2893_wire_constant & nacc1_3293_2894_buffered;
      req <= phi_stmt_2889_req_0 & phi_stmt_2889_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2889",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2889_ack_0,
          idata => idata,
          odata => acc1_2889,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2889
    phi_stmt_2895: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2898_wire_constant & nacc2_3302_2899_buffered;
      req <= phi_stmt_2895_req_0 & phi_stmt_2895_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2895",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2895_ack_0,
          idata => idata,
          odata => acc2_2895,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2895
    phi_stmt_2900: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2903_wire_constant & n_row_3284_2904_buffered;
      req <= phi_stmt_2900_req_0 & phi_stmt_2900_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2900",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2900_ack_0,
          idata => idata,
          odata => row_2900,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2900
    phi_stmt_2905: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2908_wire_constant & n_col_3276_2909_buffered;
      req <= phi_stmt_2905_req_0 & phi_stmt_2905_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2905",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2905_ack_0,
          idata => idata,
          odata => col_2905,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2905
    phi_stmt_2910: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2913_wire_constant & n_num_3265_2914_buffered;
      req <= phi_stmt_2910_req_0 & phi_stmt_2910_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2910",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2910_ack_0,
          idata => idata,
          odata => num_2910,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2910
    phi_stmt_2915: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2918_wire_constant & n_chl_3254_2919_buffered;
      req <= phi_stmt_2915_req_0 & phi_stmt_2915_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2915",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2915_ack_0,
          idata => idata,
          odata => chl_2915,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2915
    -- flow-through select operator MUX_2969_inst
    iread1_2970 <= temp2_1_2933 when (read_ip_2906_delayed_1_0_2964(0) /=  '0') else temp1_1_2949;
    -- flow-through select operator MUX_2978_inst
    iread2_2979 <= temp2_2_2937 when (read_ip_2912_delayed_1_0_2973(0) /=  '0') else temp1_2_2953;
    -- flow-through select operator MUX_2987_inst
    iread3_2988 <= temp2_3_2941 when (read_ip_2918_delayed_1_0_2982(0) /=  '0') else temp1_3_2957;
    -- flow-through select operator MUX_2996_inst
    iread4_2997 <= temp2_4_2945 when (read_ip_2924_delayed_1_0_2991(0) /=  '0') else temp1_4_2961;
    -- flow-through select operator MUX_3091_inst
    kread1_3092 <= tempk1_1_3063 when (read_k_3004_delayed_1_0_3086(0) /=  '0') else tempk2_1_3075;
    -- flow-through select operator MUX_3100_inst
    kread2_3101 <= tempk1_2_3067 when (read_k_3010_delayed_1_0_3095(0) /=  '0') else tempk2_2_3079;
    -- flow-through select operator MUX_3109_inst
    kread3_3110 <= tempk1_3_3071 when (read_k_3016_delayed_1_0_3104(0) /=  '0') else tempk2_3_3083;
    -- flow-through select operator MUX_3253_inst
    n_chl_3254 <= konst_3249_wire_constant when (chl_done_3187(0) /=  '0') else ADD_u16_u16_3252_wire;
    -- flow-through select operator MUX_3262_inst
    MUX_3262_wire <= konst_3258_wire_constant when (num_done_3194(0) /=  '0') else ADD_u2_u2_3261_wire;
    -- flow-through select operator MUX_3264_inst
    n_num_3265 <= MUX_3262_wire when (chl_done_3187(0) /=  '0') else num_2910;
    -- flow-through select operator MUX_3273_inst
    MUX_3273_wire <= konst_3269_wire_constant when (col_done_3199(0) /=  '0') else ADD_u16_u16_3272_wire;
    -- flow-through select operator MUX_3275_inst
    n_col_3276 <= MUX_3273_wire when (num_done_3194(0) /=  '0') else col_2905;
    -- flow-through select operator MUX_3283_inst
    n_row_3284 <= ADD_u16_u16_3281_wire when (row_done_3204(0) /=  '0') else row_2900;
    -- flow-through select operator MUX_3292_inst
    nacc1_3293 <= konst_3290_wire_constant when (num_done_3178_delayed_1_0_3287(0) /=  '0') else acc_val1_3170;
    -- flow-through select operator MUX_3301_inst
    nacc2_3302 <= konst_3299_wire_constant when (num_done_3184_delayed_1_0_3296(0) /=  '0') else acc_val2_3182;
    W_acc1_3070_delayed_1_0_3159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc1_3070_delayed_1_0_3159_inst_req_0;
      W_acc1_3070_delayed_1_0_3159_inst_ack_0<= wack(0);
      rreq(0) <= W_acc1_3070_delayed_1_0_3159_inst_req_1;
      W_acc1_3070_delayed_1_0_3159_inst_ack_1<= rack(0);
      W_acc1_3070_delayed_1_0_3159_inst : InterlockBuffer generic map ( -- 
        name => "W_acc1_3070_delayed_1_0_3159_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc1_2889,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc1_3070_delayed_1_0_3161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_acc2_3079_delayed_1_0_3171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc2_3079_delayed_1_0_3171_inst_req_0;
      W_acc2_3079_delayed_1_0_3171_inst_ack_0<= wack(0);
      rreq(0) <= W_acc2_3079_delayed_1_0_3171_inst_req_1;
      W_acc2_3079_delayed_1_0_3171_inst_ack_1<= rack(0);
      W_acc2_3079_delayed_1_0_3171_inst : InterlockBuffer generic map ( -- 
        name => "W_acc2_3079_delayed_1_0_3171_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc2_2895,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc2_3079_delayed_1_0_3173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_3178_delayed_1_0_3285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_3178_delayed_1_0_3285_inst_req_0;
      W_num_done_3178_delayed_1_0_3285_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_3178_delayed_1_0_3285_inst_req_1;
      W_num_done_3178_delayed_1_0_3285_inst_ack_1<= rack(0);
      W_num_done_3178_delayed_1_0_3285_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_3178_delayed_1_0_3285_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_3194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_3178_delayed_1_0_3287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_3184_delayed_1_0_3294_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_3184_delayed_1_0_3294_inst_req_0;
      W_num_done_3184_delayed_1_0_3294_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_3184_delayed_1_0_3294_inst_req_1;
      W_num_done_3184_delayed_1_0_3294_inst_ack_1<= rack(0);
      W_num_done_3184_delayed_1_0_3294_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_3184_delayed_1_0_3294_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_3194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_3184_delayed_1_0_3296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_3189_delayed_1_0_3303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_3189_delayed_1_0_3303_inst_req_0;
      W_num_done_3189_delayed_1_0_3303_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_3189_delayed_1_0_3303_inst_req_1;
      W_num_done_3189_delayed_1_0_3303_inst_ack_1<= rack(0);
      W_num_done_3189_delayed_1_0_3303_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_3189_delayed_1_0_3303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_3194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_3189_delayed_1_0_3305,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_3194_delayed_1_0_3311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_3194_delayed_1_0_3311_inst_req_0;
      W_num_done_3194_delayed_1_0_3311_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_3194_delayed_1_0_3311_inst_req_1;
      W_num_done_3194_delayed_1_0_3311_inst_ack_1<= rack(0);
      W_num_done_3194_delayed_1_0_3311_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_3194_delayed_1_0_3311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_3194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_3194_delayed_1_0_3313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2906_delayed_1_0_2962_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2906_delayed_1_0_2962_inst_req_0;
      W_read_ip_2906_delayed_1_0_2962_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2906_delayed_1_0_2962_inst_req_1;
      W_read_ip_2906_delayed_1_0_2962_inst_ack_1<= rack(0);
      W_read_ip_2906_delayed_1_0_2962_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2906_delayed_1_0_2962_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2929,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2906_delayed_1_0_2964,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2912_delayed_1_0_2971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2912_delayed_1_0_2971_inst_req_0;
      W_read_ip_2912_delayed_1_0_2971_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2912_delayed_1_0_2971_inst_req_1;
      W_read_ip_2912_delayed_1_0_2971_inst_ack_1<= rack(0);
      W_read_ip_2912_delayed_1_0_2971_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2912_delayed_1_0_2971_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2929,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2912_delayed_1_0_2973,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2918_delayed_1_0_2980_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2918_delayed_1_0_2980_inst_req_0;
      W_read_ip_2918_delayed_1_0_2980_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2918_delayed_1_0_2980_inst_req_1;
      W_read_ip_2918_delayed_1_0_2980_inst_ack_1<= rack(0);
      W_read_ip_2918_delayed_1_0_2980_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2918_delayed_1_0_2980_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2929,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2918_delayed_1_0_2982,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2924_delayed_1_0_2989_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2924_delayed_1_0_2989_inst_req_0;
      W_read_ip_2924_delayed_1_0_2989_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2924_delayed_1_0_2989_inst_req_1;
      W_read_ip_2924_delayed_1_0_2989_inst_ack_1<= rack(0);
      W_read_ip_2924_delayed_1_0_2989_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2924_delayed_1_0_2989_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2929,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2924_delayed_1_0_2991,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_3004_delayed_1_0_3084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_3004_delayed_1_0_3084_inst_req_0;
      W_read_k_3004_delayed_1_0_3084_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_3004_delayed_1_0_3084_inst_req_1;
      W_read_k_3004_delayed_1_0_3084_inst_ack_1<= rack(0);
      W_read_k_3004_delayed_1_0_3084_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_3004_delayed_1_0_3084_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_3059,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_3004_delayed_1_0_3086,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_3010_delayed_1_0_3093_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_3010_delayed_1_0_3093_inst_req_0;
      W_read_k_3010_delayed_1_0_3093_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_3010_delayed_1_0_3093_inst_req_1;
      W_read_k_3010_delayed_1_0_3093_inst_ack_1<= rack(0);
      W_read_k_3010_delayed_1_0_3093_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_3010_delayed_1_0_3093_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_3059,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_3010_delayed_1_0_3095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_3016_delayed_1_0_3102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_3016_delayed_1_0_3102_inst_req_0;
      W_read_k_3016_delayed_1_0_3102_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_3016_delayed_1_0_3102_inst_req_1;
      W_read_k_3016_delayed_1_0_3102_inst_ack_1<= rack(0);
      W_read_k_3016_delayed_1_0_3102_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_3016_delayed_1_0_3102_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_3059,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_3016_delayed_1_0_3104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_3127_delayed_1_0_3226_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_3127_delayed_1_0_3226_inst_req_0;
      W_store_kernel_3127_delayed_1_0_3226_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_3127_delayed_1_0_3226_inst_req_1;
      W_store_kernel_3127_delayed_1_0_3226_inst_ack_1<= rack(0);
      W_store_kernel_3127_delayed_1_0_3226_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_3127_delayed_1_0_3226_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_3220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_3127_delayed_1_0_3228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_3131_delayed_1_0_3233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_3131_delayed_1_0_3233_inst_req_0;
      W_store_kernel_3131_delayed_1_0_3233_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_3131_delayed_1_0_3233_inst_req_1;
      W_store_kernel_3131_delayed_1_0_3233_inst_ack_1<= rack(0);
      W_store_kernel_3131_delayed_1_0_3233_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_3131_delayed_1_0_3233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_3220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_3131_delayed_1_0_3235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_3135_delayed_1_0_3240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_3135_delayed_1_0_3240_inst_req_0;
      W_store_kernel_3135_delayed_1_0_3240_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_3135_delayed_1_0_3240_inst_req_1;
      W_store_kernel_3135_delayed_1_0_3240_inst_ack_1<= rack(0);
      W_store_kernel_3135_delayed_1_0_3240_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_3135_delayed_1_0_3240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_3220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_3135_delayed_1_0_3242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2938_delayed_1_0_3007_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2938_delayed_1_0_3007_inst_req_0;
      W_write_input_2938_delayed_1_0_3007_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2938_delayed_1_0_3007_inst_req_1;
      W_write_input_2938_delayed_1_0_3007_inst_ack_1<= rack(0);
      W_write_input_2938_delayed_1_0_3007_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2938_delayed_1_0_3007_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_3006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2938_delayed_1_0_3009,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2942_delayed_1_0_3014_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2942_delayed_1_0_3014_inst_req_0;
      W_write_input_2942_delayed_1_0_3014_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2942_delayed_1_0_3014_inst_req_1;
      W_write_input_2942_delayed_1_0_3014_inst_ack_1<= rack(0);
      W_write_input_2942_delayed_1_0_3014_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2942_delayed_1_0_3014_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_3006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2942_delayed_1_0_3016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2946_delayed_1_0_3021_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2946_delayed_1_0_3021_inst_req_0;
      W_write_input_2946_delayed_1_0_3021_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2946_delayed_1_0_3021_inst_req_1;
      W_write_input_2946_delayed_1_0_3021_inst_ack_1<= rack(0);
      W_write_input_2946_delayed_1_0_3021_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2946_delayed_1_0_3021_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_3006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2946_delayed_1_0_3023,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2950_delayed_1_0_3028_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2950_delayed_1_0_3028_inst_req_0;
      W_write_input_2950_delayed_1_0_3028_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2950_delayed_1_0_3028_inst_req_1;
      W_write_input_2950_delayed_1_0_3028_inst_ack_1<= rack(0);
      W_write_input_2950_delayed_1_0_3028_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2950_delayed_1_0_3028_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_3006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2950_delayed_1_0_3030,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_3254_2919_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_3254_2919_buf_req_0;
      n_chl_3254_2919_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_3254_2919_buf_req_1;
      n_chl_3254_2919_buf_ack_1<= rack(0);
      n_chl_3254_2919_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_3254_2919_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_3254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_3254_2919_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_3276_2909_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_3276_2909_buf_req_0;
      n_col_3276_2909_buf_ack_0<= wack(0);
      rreq(0) <= n_col_3276_2909_buf_req_1;
      n_col_3276_2909_buf_ack_1<= rack(0);
      n_col_3276_2909_buf : InterlockBuffer generic map ( -- 
        name => "n_col_3276_2909_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_3276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_3276_2909_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_num_3265_2914_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_num_3265_2914_buf_req_0;
      n_num_3265_2914_buf_ack_0<= wack(0);
      rreq(0) <= n_num_3265_2914_buf_req_1;
      n_num_3265_2914_buf_ack_1<= rack(0);
      n_num_3265_2914_buf : InterlockBuffer generic map ( -- 
        name => "n_num_3265_2914_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_num_3265,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_num_3265_2914_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_3284_2904_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_3284_2904_buf_req_0;
      n_row_3284_2904_buf_ack_0<= wack(0);
      rreq(0) <= n_row_3284_2904_buf_req_1;
      n_row_3284_2904_buf_ack_1<= rack(0);
      n_row_3284_2904_buf : InterlockBuffer generic map ( -- 
        name => "n_row_3284_2904_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_3284,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_3284_2904_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc1_3293_2894_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc1_3293_2894_buf_req_0;
      nacc1_3293_2894_buf_ack_0<= wack(0);
      rreq(0) <= nacc1_3293_2894_buf_req_1;
      nacc1_3293_2894_buf_ack_1<= rack(0);
      nacc1_3293_2894_buf : InterlockBuffer generic map ( -- 
        name => "nacc1_3293_2894_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc1_3293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc1_3293_2894_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc2_3302_2899_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc2_3302_2899_buf_req_0;
      nacc2_3302_2899_buf_ack_0<= wack(0);
      rreq(0) <= nacc2_3302_2899_buf_req_1;
      nacc2_3302_2899_buf_ack_1<= rack(0);
      nacc2_3302_2899_buf : InterlockBuffer generic map ( -- 
        name => "nacc2_3302_2899_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc2_3302,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc2_3302_2899_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3037_inst
    process(iread1_2970) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread1_2970(15 downto 0);
      ival1_3038 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3041_inst
    process(iread2_2979) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread2_2979(15 downto 0);
      ival2_3042 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3045_inst
    process(iread3_2988) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread3_2988(15 downto 0);
      ival3_3046 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3049_inst
    process(iread4_2997) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread4_2997(15 downto 0);
      ival4_3050 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3113_inst
    process(kread1_3092) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread1_3092(15 downto 0);
      kval1_3114 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3117_inst
    process(kread2_3101) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread2_3101(15 downto 0);
      kval2_3118 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3121_inst
    process(kread3_3110) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread3_3110(15 downto 0);
      kval3_3122 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3127_inst
    process(MUL_i16_i16_3126_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_3126_wire(15 downto 0);
      mul_val1_3128 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3133_inst
    process(MUL_i16_i16_3132_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_3132_wire(15 downto 0);
      mul_val2_3134 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3139_inst
    process(MUL_i16_i16_3138_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_3138_wire(15 downto 0);
      mul_val3_3140 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3145_inst
    process(MUL_i16_i16_3144_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_3144_wire(15 downto 0);
      mul_val4_3146 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3151_inst
    process(MUL_i16_i16_3150_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_3150_wire(15 downto 0);
      mul_val5_3152 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3157_inst
    process(MUL_i16_i16_3156_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_3156_wire(15 downto 0);
      mul_val6_3158 <= tmp_var; -- 
    end process;
    type_cast_3309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_3309_inst_req_0;
      type_cast_3309_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_3309_inst_req_1;
      type_cast_3309_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  num_done_3189_delayed_1_0_3305(0);
      type_cast_3309_inst_gI: SplitGuardInterface generic map(name => "type_cast_3309_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_3309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val1_3170,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3309_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3317_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_3317_inst_req_0;
      type_cast_3317_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_3317_inst_req_1;
      type_cast_3317_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  num_done_3194_delayed_1_0_3313(0);
      type_cast_3317_inst_gI: SplitGuardInterface generic map(name => "type_cast_3317_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_3317_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3317_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val2_3182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3317_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_2887_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_3321_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2887_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2887_branch_req_0,
          ack0 => do_while_stmt_2887_branch_ack_0,
          ack1 => do_while_stmt_2887_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_3165_inst
    process(acc1_3070_delayed_1_0_3161, mul_val1_3128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc1_3070_delayed_1_0_3161, mul_val1_3128, tmp_var);
      ADD_i16_i16_3165_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_3168_inst
    process(mul_val2_3134, mul_val3_3140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val2_3134, mul_val3_3140, tmp_var);
      ADD_i16_i16_3168_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_3169_inst
    process(ADD_i16_i16_3165_wire, ADD_i16_i16_3168_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i16_i16_3165_wire, ADD_i16_i16_3168_wire, tmp_var);
      acc_val1_3170 <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_3177_inst
    process(acc2_3079_delayed_1_0_3173, mul_val4_3146) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc2_3079_delayed_1_0_3173, mul_val4_3146, tmp_var);
      ADD_i16_i16_3177_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_3180_inst
    process(mul_val5_3152, mul_val6_3158) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_3152, mul_val6_3158, tmp_var);
      ADD_i16_i16_3180_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_3181_inst
    process(ADD_i16_i16_3177_wire, ADD_i16_i16_3180_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i16_i16_3177_wire, ADD_i16_i16_3180_wire, tmp_var);
      acc_val2_3182 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3252_inst
    process(chl_2915) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_2915, konst_3251_wire_constant, tmp_var);
      ADD_u16_u16_3252_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3272_inst
    process(col_2905) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_2905, konst_3271_wire_constant, tmp_var);
      ADD_u16_u16_3272_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3281_inst
    process(row_2900) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_2900, konst_3280_wire_constant, tmp_var);
      ADD_u16_u16_3281_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u2_u2_3261_inst
    process(num_2910) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_2910, konst_3260_wire_constant, tmp_var);
      ADD_u2_u2_3261_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3005_inst
    process(ULT_u16_u1_3001_wire, UGT_u2_u1_3004_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ULT_u16_u1_3001_wire, UGT_u2_u1_3004_wire, tmp_var);
      write_input_3006 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3058_inst
    process(EQ_u16_u1_3054_wire, EQ_u16_u1_3057_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u16_u1_3054_wire, EQ_u16_u1_3057_wire, tmp_var);
      read_k_3059 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3193_inst
    process(EQ_u2_u1_3191_wire, chl_done_3187) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_3191_wire, chl_done_3187, tmp_var);
      num_done_3194 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3203_inst
    process(col_done_3199, num_done_3194) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_3199, num_done_3194, tmp_var);
      row_done_3204 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3218_inst
    process(out_done_flag_3214, col_done_3199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_3214, col_done_3199, tmp_var);
      AND_u1_u1_3218_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3224_inst
    process(out_done_flag_3214, row_done_3204) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_3214, row_done_3204, tmp_var);
      all_done_flag_3225 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2924_inst
    process(col_2905) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2905, konst_2923_wire_constant, tmp_var);
      EQ_u16_u1_2924_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_3054_inst
    process(col_2905) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2905, konst_3053_wire_constant, tmp_var);
      EQ_u16_u1_3054_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_3057_inst
    process(row_2900) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(row_2900, konst_3056_wire_constant, tmp_var);
      EQ_u16_u1_3057_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_3186_inst
    process(chl_2915, num_chl_2886) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(chl_2915, num_chl_2886, tmp_var);
      chl_done_3187 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_3198_inst
    process(col_2905, num_col_2881) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2905, num_col_2881, tmp_var);
      col_done_3199 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2927_inst
    process(num_2910) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_2910, konst_2926_wire_constant, tmp_var);
      EQ_u2_u1_2927_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_3191_inst
    process(num_2910) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_2910, konst_3190_wire_constant, tmp_var);
      EQ_u2_u1_3191_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_3126_inst
    process(kval1_3114, ival1_3038) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_3114, ival1_3038, tmp_var);
      MUL_i16_i16_3126_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_3132_inst
    process(kval2_3118, ival2_3042) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_3118, ival2_3042, tmp_var);
      MUL_i16_i16_3132_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_3138_inst
    process(kval3_3122, ival3_3046) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_3122, ival3_3046, tmp_var);
      MUL_i16_i16_3138_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_3144_inst
    process(kval1_3114, ival2_3042) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_3114, ival2_3042, tmp_var);
      MUL_i16_i16_3144_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_3150_inst
    process(kval2_3118, ival3_3046) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_3118, ival3_3046, tmp_var);
      MUL_i16_i16_3150_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_3156_inst
    process(kval3_3122, ival4_3050) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_3122, ival4_3050, tmp_var);
      MUL_i16_i16_3156_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_3219_inst
    process(AND_u1_u1_3218_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AND_u1_u1_3218_wire, tmp_var);
      store_kernel_3220 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3321_inst
    process(all_done_flag_3225) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", all_done_flag_3225, tmp_var);
      NOT_u1_u1_3321_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2928_inst
    process(EQ_u16_u1_2924_wire, EQ_u2_u1_2927_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u16_u1_2924_wire, EQ_u2_u1_2927_wire, tmp_var);
      read_ip_2929 <= tmp_var; --
    end process;
    -- shared split operator group (32) : SUB_u16_u16_2875_inst 
    ApIntSub_group_32: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_2873_wire;
      num_row_2876 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2875_inst_req_0;
      SUB_u16_u16_2875_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2875_inst_req_1;
      SUB_u16_u16_2875_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_32_gI: SplitGuardInterface generic map(name => "ApIntSub_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : SUB_u16_u16_2880_inst 
    ApIntSub_group_33: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_2878_wire;
      num_col_2881 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2880_inst_req_0;
      SUB_u16_u16_2880_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2880_inst_req_1;
      SUB_u16_u16_2880_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_33_gI: SplitGuardInterface generic map(name => "ApIntSub_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : SUB_u16_u16_2885_inst 
    ApIntSub_group_34: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_size_pipe_2883_wire;
      num_chl_2886 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2885_inst_req_0;
      SUB_u16_u16_2885_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2885_inst_req_1;
      SUB_u16_u16_2885_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_34_gI: SplitGuardInterface generic map(name => "ApIntSub_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : SUB_u16_u16_3208_inst 
    ApIntSub_group_35: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= num_row_2876;
      SUB_u16_u16_3113_3113_delayed_1_0_3209 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3208_inst_req_0;
      SUB_u16_u16_3208_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3208_inst_req_1;
      SUB_u16_u16_3208_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_35_gI: SplitGuardInterface generic map(name => "ApIntSub_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- binary operator UGE_u16_u1_3213_inst
    process(row_2900, SUB_u16_u16_3113_3113_delayed_1_0_3209) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(row_2900, SUB_u16_u16_3113_3113_delayed_1_0_3209, tmp_var);
      out_done_flag_3214 <= tmp_var; --
    end process;
    -- binary operator UGT_u2_u1_3004_inst
    process(num_2910) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_2910, konst_3003_wire_constant, tmp_var);
      UGT_u2_u1_3004_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_3001_inst
    process(col_2905, num_col_2881) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(col_2905, num_col_2881, tmp_var);
      ULT_u16_u1_3001_wire <= tmp_var; --
    end process;
    xxconvolvexxconv_ip1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip1",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip1_pipe_read_req,
        read_ack => xxconvolvexxconv_ip1_pipe_read_ack,
        read_data => xxconvolvexxconv_ip1_pipe_read_data,
        write_req => xxconvolvexxconv_ip1_pipe_write_req,
        write_ack => xxconvolvexxconv_ip1_pipe_write_ack,
        write_data => xxconvolvexxconv_ip1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip2",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip2_pipe_read_req,
        read_ack => xxconvolvexxconv_ip2_pipe_read_ack,
        read_data => xxconvolvexxconv_ip2_pipe_read_data,
        write_req => xxconvolvexxconv_ip2_pipe_write_req,
        write_ack => xxconvolvexxconv_ip2_pipe_write_ack,
        write_data => xxconvolvexxconv_ip2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip3",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip3_pipe_read_req,
        read_ack => xxconvolvexxconv_ip3_pipe_read_ack,
        read_data => xxconvolvexxconv_ip3_pipe_read_data,
        write_req => xxconvolvexxconv_ip3_pipe_write_req,
        write_ack => xxconvolvexxconv_ip3_pipe_write_ack,
        write_data => xxconvolvexxconv_ip3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip4_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip4",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip4_pipe_read_req,
        read_ack => xxconvolvexxconv_ip4_pipe_read_ack,
        read_data => xxconvolvexxconv_ip4_pipe_read_data,
        write_req => xxconvolvexxconv_ip4_pipe_write_req,
        write_ack => xxconvolvexxconv_ip4_pipe_write_ack,
        write_data => xxconvolvexxconv_ip4_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k1",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k1_pipe_read_req,
        read_ack => xxconvolvexxconv_k1_pipe_read_ack,
        read_data => xxconvolvexxconv_k1_pipe_read_data,
        write_req => xxconvolvexxconv_k1_pipe_write_req,
        write_ack => xxconvolvexxconv_k1_pipe_write_ack,
        write_data => xxconvolvexxconv_k1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k2",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k2_pipe_read_req,
        read_ack => xxconvolvexxconv_k2_pipe_read_ack,
        read_data => xxconvolvexxconv_k2_pipe_read_data,
        write_req => xxconvolvexxconv_k2_pipe_write_req,
        write_ack => xxconvolvexxconv_k2_pipe_write_ack,
        write_data => xxconvolvexxconv_k2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k3",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k3_pipe_read_req,
        read_ack => xxconvolvexxconv_k3_pipe_read_ack,
        read_data => xxconvolvexxconv_k3_pipe_read_data,
        write_req => xxconvolvexxconv_k3_pipe_write_req,
        write_ack => xxconvolvexxconv_k3_pipe_write_ack,
        write_data => xxconvolvexxconv_k3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : RPIPE_input_pipe1_2932_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_2932_inst_req_0;
      RPIPE_input_pipe1_2932_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_2932_inst_req_1;
      RPIPE_input_pipe1_2932_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2929(0);
      temp2_1_2933 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_input_pipe2_2936_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe2_2936_inst_req_0;
      RPIPE_input_pipe2_2936_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe2_2936_inst_req_1;
      RPIPE_input_pipe2_2936_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2929(0);
      temp2_2_2937 <= data_out(15 downto 0);
      input_pipe2_read_1_gI: SplitGuardInterface generic map(name => "input_pipe2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe2_read_1: InputPortRevised -- 
        generic map ( name => "input_pipe2_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe2_pipe_read_req(0),
          oack => input_pipe2_pipe_read_ack(0),
          odata => input_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_input_pipe3_2940_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe3_2940_inst_req_0;
      RPIPE_input_pipe3_2940_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe3_2940_inst_req_1;
      RPIPE_input_pipe3_2940_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2929(0);
      temp2_3_2941 <= data_out(15 downto 0);
      input_pipe3_read_2_gI: SplitGuardInterface generic map(name => "input_pipe3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe3_read_2: InputPortRevised -- 
        generic map ( name => "input_pipe3_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe3_pipe_read_req(0),
          oack => input_pipe3_pipe_read_ack(0),
          odata => input_pipe3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_input_pipe4_2944_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe4_2944_inst_req_0;
      RPIPE_input_pipe4_2944_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe4_2944_inst_req_1;
      RPIPE_input_pipe4_2944_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2929(0);
      temp2_4_2945 <= data_out(15 downto 0);
      input_pipe4_read_3_gI: SplitGuardInterface generic map(name => "input_pipe4_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe4_read_3: InputPortRevised -- 
        generic map ( name => "input_pipe4_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe4_pipe_read_req(0),
          oack => input_pipe4_pipe_read_ack(0),
          odata => input_pipe4_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_kernel_pipe1_3062_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_3062_inst_req_0;
      RPIPE_kernel_pipe1_3062_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_3062_inst_req_1;
      RPIPE_kernel_pipe1_3062_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_3059(0);
      tempk1_1_3063 <= data_out(15 downto 0);
      kernel_pipe1_read_4_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_4: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_4", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : RPIPE_kernel_pipe2_3066_inst 
    InportGroup_5: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe2_3066_inst_req_0;
      RPIPE_kernel_pipe2_3066_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe2_3066_inst_req_1;
      RPIPE_kernel_pipe2_3066_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_3059(0);
      tempk1_2_3067 <= data_out(15 downto 0);
      kernel_pipe2_read_5_gI: SplitGuardInterface generic map(name => "kernel_pipe2_read_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_read_5: InputPortRevised -- 
        generic map ( name => "kernel_pipe2_read_5", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe2_pipe_read_req(0),
          oack => kernel_pipe2_pipe_read_ack(0),
          odata => kernel_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : RPIPE_kernel_pipe3_3070_inst 
    InportGroup_6: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe3_3070_inst_req_0;
      RPIPE_kernel_pipe3_3070_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe3_3070_inst_req_1;
      RPIPE_kernel_pipe3_3070_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_3059(0);
      tempk1_3_3071 <= data_out(15 downto 0);
      kernel_pipe3_read_6_gI: SplitGuardInterface generic map(name => "kernel_pipe3_read_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_read_6: InputPortRevised -- 
        generic map ( name => "kernel_pipe3_read_6", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe3_pipe_read_req(0),
          oack => kernel_pipe3_pipe_read_ack(0),
          odata => kernel_pipe3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : RPIPE_num_out_pipe_2878_inst RPIPE_num_out_pipe_2873_inst 
    InportGroup_7: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_num_out_pipe_2878_inst_req_0;
      reqL_unguarded(0) <= RPIPE_num_out_pipe_2873_inst_req_0;
      RPIPE_num_out_pipe_2878_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_num_out_pipe_2873_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_num_out_pipe_2878_inst_req_1;
      reqR_unguarded(0) <= RPIPE_num_out_pipe_2873_inst_req_1;
      RPIPE_num_out_pipe_2878_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_num_out_pipe_2873_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      RPIPE_num_out_pipe_2878_wire <= data_out(31 downto 16);
      RPIPE_num_out_pipe_2873_wire <= data_out(15 downto 0);
      num_out_pipe_read_7_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_7_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_7: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_7", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : RPIPE_size_pipe_2883_inst 
    InportGroup_8: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_2883_inst_req_0;
      RPIPE_size_pipe_2883_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_2883_inst_req_1;
      RPIPE_size_pipe_2883_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_size_pipe_2883_wire <= data_out(15 downto 0);
      size_pipe_read_8_gI: SplitGuardInterface generic map(name => "size_pipe_read_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_8: InputPortRevised -- 
        generic map ( name => "size_pipe_read_8", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : RPIPE_xxconvolvexxconv_ip1_2948_inst 
    InportGroup_9: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_2948_inst_req_0;
      RPIPE_xxconvolvexxconv_ip1_2948_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_2948_inst_req_1;
      RPIPE_xxconvolvexxconv_ip1_2948_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2929(0);
      temp1_1_2949 <= data_out(15 downto 0);
      xxconvolvexxconv_ip1_read_9_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_read_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_read_9: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1_read_9", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip1_pipe_read_req(0),
          oack => xxconvolvexxconv_ip1_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : RPIPE_xxconvolvexxconv_ip2_2952_inst 
    InportGroup_10: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_2952_inst_req_0;
      RPIPE_xxconvolvexxconv_ip2_2952_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_2952_inst_req_1;
      RPIPE_xxconvolvexxconv_ip2_2952_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2929(0);
      temp1_2_2953 <= data_out(15 downto 0);
      xxconvolvexxconv_ip2_read_10_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_read_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_read_10: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2_read_10", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip2_pipe_read_req(0),
          oack => xxconvolvexxconv_ip2_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : RPIPE_xxconvolvexxconv_ip3_2956_inst 
    InportGroup_11: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_2956_inst_req_0;
      RPIPE_xxconvolvexxconv_ip3_2956_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_2956_inst_req_1;
      RPIPE_xxconvolvexxconv_ip3_2956_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2929(0);
      temp1_3_2957 <= data_out(15 downto 0);
      xxconvolvexxconv_ip3_read_11_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_read_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_read_11: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3_read_11", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip3_pipe_read_req(0),
          oack => xxconvolvexxconv_ip3_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- shared inport operator group (12) : RPIPE_xxconvolvexxconv_ip4_2960_inst 
    InportGroup_12: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip4_2960_inst_req_0;
      RPIPE_xxconvolvexxconv_ip4_2960_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip4_2960_inst_req_1;
      RPIPE_xxconvolvexxconv_ip4_2960_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2929(0);
      temp1_4_2961 <= data_out(15 downto 0);
      xxconvolvexxconv_ip4_read_12_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip4_read_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip4_read_12: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip4_read_12", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip4_pipe_read_req(0),
          oack => xxconvolvexxconv_ip4_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip4_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 12
    -- shared inport operator group (13) : RPIPE_xxconvolvexxconv_k1_3074_inst 
    InportGroup_13: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_3074_inst_req_0;
      RPIPE_xxconvolvexxconv_k1_3074_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_3074_inst_req_1;
      RPIPE_xxconvolvexxconv_k1_3074_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_3059(0);
      tempk2_1_3075 <= data_out(15 downto 0);
      xxconvolvexxconv_k1_read_13_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_read_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_read_13: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1_read_13", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k1_pipe_read_req(0),
          oack => xxconvolvexxconv_k1_pipe_read_ack(0),
          odata => xxconvolvexxconv_k1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 13
    -- shared inport operator group (14) : RPIPE_xxconvolvexxconv_k2_3078_inst 
    InportGroup_14: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_3078_inst_req_0;
      RPIPE_xxconvolvexxconv_k2_3078_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_3078_inst_req_1;
      RPIPE_xxconvolvexxconv_k2_3078_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_3059(0);
      tempk2_2_3079 <= data_out(15 downto 0);
      xxconvolvexxconv_k2_read_14_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_read_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_read_14: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2_read_14", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k2_pipe_read_req(0),
          oack => xxconvolvexxconv_k2_pipe_read_ack(0),
          odata => xxconvolvexxconv_k2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 14
    -- shared inport operator group (15) : RPIPE_xxconvolvexxconv_k3_3082_inst 
    InportGroup_15: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_3082_inst_req_0;
      RPIPE_xxconvolvexxconv_k3_3082_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_3082_inst_req_1;
      RPIPE_xxconvolvexxconv_k3_3082_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_3059(0);
      tempk2_3_3083 <= data_out(15 downto 0);
      xxconvolvexxconv_k3_read_15_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_read_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_read_15: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3_read_15", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k3_pipe_read_req(0),
          oack => xxconvolvexxconv_k3_pipe_read_ack(0),
          odata => xxconvolvexxconv_k3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 15
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3322_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3322_inst_req_0;
      WPIPE_input_done_pipe_3322_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3322_inst_req_1;
      WPIPE_input_done_pipe_3322_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3323_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_output_pipe_3307_inst WPIPE_output_pipe_3315_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_output_pipe_3307_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_output_pipe_3315_inst_req_0;
      WPIPE_output_pipe_3307_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_output_pipe_3315_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_output_pipe_3307_inst_req_1;
      update_req_unguarded(0) <= WPIPE_output_pipe_3315_inst_req_1;
      WPIPE_output_pipe_3307_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_output_pipe_3315_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= num_done_3194_delayed_1_0_3313(0);
      guard_vector(1)  <= num_done_3189_delayed_1_0_3305(0);
      data_in <= type_cast_3309_wire & type_cast_3317_wire;
      output_pipe_write_1_gI: SplitGuardInterface generic map(name => "output_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_xxconvolvexxconv_ip1_3011_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_3011_inst_req_0;
      WPIPE_xxconvolvexxconv_ip1_3011_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_3011_inst_req_1;
      WPIPE_xxconvolvexxconv_ip1_3011_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2938_delayed_1_0_3009(0);
      data_in <= iread1_2970;
      xxconvolvexxconv_ip1_write_2_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_write_2: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip1_pipe_write_req(0),
          oack => xxconvolvexxconv_ip1_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_xxconvolvexxconv_ip2_3018_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_3018_inst_req_0;
      WPIPE_xxconvolvexxconv_ip2_3018_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_3018_inst_req_1;
      WPIPE_xxconvolvexxconv_ip2_3018_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2942_delayed_1_0_3016(0);
      data_in <= iread2_2979;
      xxconvolvexxconv_ip2_write_3_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_write_3: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip2_pipe_write_req(0),
          oack => xxconvolvexxconv_ip2_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_xxconvolvexxconv_ip3_3025_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_3025_inst_req_0;
      WPIPE_xxconvolvexxconv_ip3_3025_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_3025_inst_req_1;
      WPIPE_xxconvolvexxconv_ip3_3025_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2946_delayed_1_0_3023(0);
      data_in <= iread3_2988;
      xxconvolvexxconv_ip3_write_4_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_write_4: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip3_pipe_write_req(0),
          oack => xxconvolvexxconv_ip3_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_xxconvolvexxconv_ip4_3032_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip4_3032_inst_req_0;
      WPIPE_xxconvolvexxconv_ip4_3032_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip4_3032_inst_req_1;
      WPIPE_xxconvolvexxconv_ip4_3032_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2950_delayed_1_0_3030(0);
      data_in <= iread4_2997;
      xxconvolvexxconv_ip4_write_5_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip4_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip4_write_5: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip4", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip4_pipe_write_req(0),
          oack => xxconvolvexxconv_ip4_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip4_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_xxconvolvexxconv_k1_3230_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_3230_inst_req_0;
      WPIPE_xxconvolvexxconv_k1_3230_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_3230_inst_req_1;
      WPIPE_xxconvolvexxconv_k1_3230_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_3127_delayed_1_0_3228(0);
      data_in <= kread1_3092;
      xxconvolvexxconv_k1_write_6_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_write_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_write_6: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k1_pipe_write_req(0),
          oack => xxconvolvexxconv_k1_pipe_write_ack(0),
          odata => xxconvolvexxconv_k1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_xxconvolvexxconv_k2_3237_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_3237_inst_req_0;
      WPIPE_xxconvolvexxconv_k2_3237_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_3237_inst_req_1;
      WPIPE_xxconvolvexxconv_k2_3237_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_3131_delayed_1_0_3235(0);
      data_in <= kread2_3101;
      xxconvolvexxconv_k2_write_7_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_write_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_write_7: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k2_pipe_write_req(0),
          oack => xxconvolvexxconv_k2_pipe_write_ack(0),
          odata => xxconvolvexxconv_k2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- shared outport operator group (8) : WPIPE_xxconvolvexxconv_k3_3244_inst 
    OutportGroup_8: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_3244_inst_req_0;
      WPIPE_xxconvolvexxconv_k3_3244_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_3244_inst_req_1;
      WPIPE_xxconvolvexxconv_k3_3244_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_3135_delayed_1_0_3242(0);
      data_in <= kread3_3110;
      xxconvolvexxconv_k3_write_8_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_write_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_write_8: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k3_pipe_write_req(0),
          oack => xxconvolvexxconv_k3_pipe_write_ack(0),
          odata => xxconvolvexxconv_k3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    num_chl : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal num_chl_buffer :  std_logic_vector(15 downto 0);
  signal num_chl_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_1909_start: Boolean;
  signal loadKernelChannel_CP_1909_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal addr_of_856_final_reg_ack_1 : boolean;
  signal ptr_deref_860_load_0_req_1 : boolean;
  signal array_obj_ref_855_index_offset_req_1 : boolean;
  signal nmycount_916_896_buf_ack_1 : boolean;
  signal addr_of_856_final_reg_ack_0 : boolean;
  signal nmycount_916_896_buf_ack_0 : boolean;
  signal ptr_deref_860_load_0_ack_0 : boolean;
  signal ptr_deref_860_load_0_req_0 : boolean;
  signal RPIPE_input_done_pipe_889_inst_req_0 : boolean;
  signal phi_stmt_894_req_0 : boolean;
  signal array_obj_ref_855_index_offset_ack_0 : boolean;
  signal do_while_stmt_892_branch_req_0 : boolean;
  signal phi_stmt_894_req_1 : boolean;
  signal phi_stmt_894_ack_0 : boolean;
  signal nmycount_916_896_buf_req_1 : boolean;
  signal RPIPE_input_done_pipe_889_inst_ack_0 : boolean;
  signal ptr_deref_860_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_889_inst_req_1 : boolean;
  signal start_add_897_buf_req_1 : boolean;
  signal array_obj_ref_855_index_offset_req_0 : boolean;
  signal addr_of_856_final_reg_req_1 : boolean;
  signal nmycount_916_896_buf_req_0 : boolean;
  signal RPIPE_input_done_pipe_889_inst_ack_1 : boolean;
  signal addr_of_856_final_reg_req_0 : boolean;
  signal start_add_897_buf_ack_0 : boolean;
  signal start_add_897_buf_req_0 : boolean;
  signal array_obj_ref_855_index_offset_ack_1 : boolean;
  signal start_add_897_buf_ack_1 : boolean;
  signal phi_stmt_898_req_1 : boolean;
  signal phi_stmt_898_req_0 : boolean;
  signal phi_stmt_898_ack_0 : boolean;
  signal my_fetch_861_900_buf_req_0 : boolean;
  signal my_fetch_861_900_buf_ack_0 : boolean;
  signal my_fetch_861_900_buf_req_1 : boolean;
  signal my_fetch_861_900_buf_ack_1 : boolean;
  signal nfetch_val_988_901_buf_req_0 : boolean;
  signal nfetch_val_988_901_buf_ack_0 : boolean;
  signal nfetch_val_988_901_buf_req_1 : boolean;
  signal nfetch_val_988_901_buf_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_942_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_942_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_942_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_942_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe2_946_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_946_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_946_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe2_946_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe3_950_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe3_950_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe3_950_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe3_950_inst_ack_1 : boolean;
  signal array_obj_ref_966_index_offset_req_0 : boolean;
  signal array_obj_ref_966_index_offset_ack_0 : boolean;
  signal array_obj_ref_966_index_offset_req_1 : boolean;
  signal array_obj_ref_966_index_offset_ack_1 : boolean;
  signal addr_of_967_final_reg_req_0 : boolean;
  signal addr_of_967_final_reg_ack_0 : boolean;
  signal addr_of_967_final_reg_req_1 : boolean;
  signal addr_of_967_final_reg_ack_1 : boolean;
  signal W_fn_921_delayed_7_0_969_inst_req_0 : boolean;
  signal W_fn_921_delayed_7_0_969_inst_ack_0 : boolean;
  signal W_fn_921_delayed_7_0_969_inst_req_1 : boolean;
  signal W_fn_921_delayed_7_0_969_inst_ack_1 : boolean;
  signal ptr_deref_975_load_0_req_0 : boolean;
  signal ptr_deref_975_load_0_ack_0 : boolean;
  signal ptr_deref_975_load_0_req_1 : boolean;
  signal ptr_deref_975_load_0_ack_1 : boolean;
  signal W_fn_927_delayed_13_0_977_inst_req_0 : boolean;
  signal W_fn_927_delayed_13_0_977_inst_ack_0 : boolean;
  signal W_fn_927_delayed_13_0_977_inst_req_1 : boolean;
  signal W_fn_927_delayed_13_0_977_inst_ack_1 : boolean;
  signal W_fetch_val_929_delayed_13_0_980_inst_req_0 : boolean;
  signal W_fetch_val_929_delayed_13_0_980_inst_ack_0 : boolean;
  signal W_fetch_val_929_delayed_13_0_980_inst_req_1 : boolean;
  signal W_fetch_val_929_delayed_13_0_980_inst_ack_1 : boolean;
  signal do_while_stmt_892_branch_ack_0 : boolean;
  signal do_while_stmt_892_branch_ack_1 : boolean;
  signal WPIPE_size_pipe_996_inst_req_0 : boolean;
  signal WPIPE_size_pipe_996_inst_ack_0 : boolean;
  signal WPIPE_size_pipe_996_inst_req_1 : boolean;
  signal WPIPE_size_pipe_996_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(79 downto 64) <= num_chl;
  num_chl_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_1909_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1909_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1909_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1909_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_1909: Block -- control-path 
    signal loadKernelChannel_CP_1909_elements: BooleanArray(98 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_1909_elements(0) <= loadKernelChannel_CP_1909_start;
    loadKernelChannel_CP_1909_symbol <= loadKernelChannel_CP_1909_elements(98);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_resized_1
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_computed_1
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_Sample/rr
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_complete/req
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_complete/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_update_start_
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_sample_start_
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_update_start_
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/$entry
      -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(0), ack => array_obj_ref_855_index_offset_req_0); -- 
    req_1959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(0), ack => addr_of_856_final_reg_req_1); -- 
    req_1944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(0), ack => array_obj_ref_855_index_offset_req_1); -- 
    cr_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(0), ack => ptr_deref_860_load_0_req_1); -- 
    rr_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(0), ack => RPIPE_input_done_pipe_889_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_Sample/ack
      -- CP-element group 1: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_Sample/$exit
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_855_index_offset_ack_0, ack => loadKernelChannel_CP_1909_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_offset_calculated
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_request/$entry
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_request/req
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_sample_start_
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_845_to_assign_stmt_890/array_obj_ref_855_final_index_sum_regn_Update/ack
      -- 
    ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_855_index_offset_ack_1, ack => loadKernelChannel_CP_1909_elements(2)); -- 
    req_1954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(2), ack => addr_of_856_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_request/ack
      -- CP-element group 3: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_sample_completed_
      -- CP-element group 3: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_request/$exit
      -- 
    ack_1955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_856_final_reg_ack_0, ack => loadKernelChannel_CP_1909_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_complete/ack
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_complete/$exit
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Sample/word_access_start/word_0/rr
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_address_resized
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/addr_of_856_update_completed_
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_sample_start_
      -- 
    ack_1960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_856_final_reg_ack_1, ack => loadKernelChannel_CP_1909_elements(4)); -- 
    rr_1993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(4), ack => ptr_deref_860_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_sample_completed_
      -- CP-element group 5: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Sample/word_access_start/$exit
      -- 
    ra_1994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_0_ack_0, ack => loadKernelChannel_CP_1909_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/$exit
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_update_completed_
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/ptr_deref_860_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/ptr_deref_860_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/ptr_deref_860_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/ptr_deref_860_Merge/merge_ack
      -- CP-element group 6: 	 assign_stmt_845_to_assign_stmt_890/ptr_deref_860_Update/word_access_complete/$exit
      -- 
    ca_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_0_ack_1, ack => loadKernelChannel_CP_1909_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_Update/$entry
      -- CP-element group 7: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_update_start_
      -- CP-element group 7: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_Sample/ra
      -- CP-element group 7: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_Update/cr
      -- CP-element group 7: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_sample_completed_
      -- 
    ra_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_889_inst_ack_0, ack => loadKernelChannel_CP_1909_elements(7)); -- 
    cr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(7), ack => RPIPE_input_done_pipe_889_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_update_completed_
      -- CP-element group 8: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_Update/$exit
      -- CP-element group 8: 	 assign_stmt_845_to_assign_stmt_890/RPIPE_input_done_pipe_889_Update/ca
      -- 
    ca_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_889_inst_ack_1, ack => loadKernelChannel_CP_1909_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_891/$entry
      -- CP-element group 9: 	 assign_stmt_845_to_assign_stmt_890/$exit
      -- CP-element group 9: 	 branch_block_stmt_891/branch_block_stmt_891__entry__
      -- CP-element group 9: 	 branch_block_stmt_891/do_while_stmt_892__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(1) & loadKernelChannel_CP_1909_elements(6) & loadKernelChannel_CP_1909_elements(8);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	96 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	97 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_891/$exit
      -- CP-element group 10: 	 branch_block_stmt_891/branch_block_stmt_891__exit__
      -- CP-element group 10: 	 branch_block_stmt_891/do_while_stmt_892__exit__
      -- CP-element group 10: 	 assign_stmt_998/$entry
      -- CP-element group 10: 	 assign_stmt_998/WPIPE_size_pipe_996_sample_start_
      -- CP-element group 10: 	 assign_stmt_998/WPIPE_size_pipe_996_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_998/WPIPE_size_pipe_996_Sample/req
      -- 
    req_2360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(10), ack => WPIPE_size_pipe_996_inst_req_0); -- 
    loadKernelChannel_CP_1909_elements(10) <= loadKernelChannel_CP_1909_elements(96);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_891/do_while_stmt_892/$entry
      -- CP-element group 11: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892__entry__
      -- 
    loadKernelChannel_CP_1909_elements(11) <= loadKernelChannel_CP_1909_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	96 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892__exit__
      -- 
    -- Element group loadKernelChannel_CP_1909_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_891/do_while_stmt_892/loop_back
      -- 
    -- Element group loadKernelChannel_CP_1909_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	94 
    -- CP-element group 14: 	95 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_891/do_while_stmt_892/condition_done
      -- CP-element group 14: 	 branch_block_stmt_891/do_while_stmt_892/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_891/do_while_stmt_892/loop_taken/$entry
      -- 
    loadKernelChannel_CP_1909_elements(14) <= loadKernelChannel_CP_1909_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	93 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_891/do_while_stmt_892/loop_body_done
      -- 
    loadKernelChannel_CP_1909_elements(15) <= loadKernelChannel_CP_1909_elements(93);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	28 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_1909_elements(16) <= loadKernelChannel_CP_1909_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_1909_elements(17) <= loadKernelChannel_CP_1909_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	70 
    -- CP-element group 18: 	71 
    -- CP-element group 18: 	92 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	42 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/loop_body_start
      -- CP-element group 18: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/$entry
      -- 
    -- Element group loadKernelChannel_CP_1909_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	92 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	27 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/condition_evaluated
      -- 
    condition_evaluated_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(19), ack => do_while_stmt_892_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(92) & loadKernelChannel_CP_1909_elements(23) & loadKernelChannel_CP_1909_elements(27);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	41 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/aggregated_phi_sample_req
      -- CP-element group 20: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_sample_start__ps
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(24) & loadKernelChannel_CP_1909_elements(41) & loadKernelChannel_CP_1909_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	81 
    -- CP-element group 21: 	85 
    -- CP-element group 21: 	89 
    -- CP-element group 21: 	93 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	41 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(26) & loadKernelChannel_CP_1909_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	42 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/aggregated_phi_update_req
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(25) & loadKernelChannel_CP_1909_elements(42);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(27) & loadKernelChannel_CP_1909_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(18) & loadKernelChannel_CP_1909_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	64 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	78 
    -- CP-element group 25: 	86 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(18) & loadKernelChannel_CP_1909_elements(61) & loadKernelChannel_CP_1909_elements(64) & loadKernelChannel_CP_1909_elements(67) & loadKernelChannel_CP_1909_elements(72) & loadKernelChannel_CP_1909_elements(78) & loadKernelChannel_CP_1909_elements(86) & loadKernelChannel_CP_1909_elements(27);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1909_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	60 
    -- CP-element group 27: 	63 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	72 
    -- CP-element group 27: 	76 
    -- CP-element group 27: 	84 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	23 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (15) 
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_resize_1/index_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_Sample/req
      -- 
    req_2226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(27), ack => array_obj_ref_966_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_1909_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	16 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_loopback_trigger
      -- 
    loadKernelChannel_CP_1909_elements(28) <= loadKernelChannel_CP_1909_elements(16);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_loopback_sample_req
      -- CP-element group 29: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_loopback_sample_req_ps
      -- 
    phi_stmt_894_loopback_sample_req_2061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_894_loopback_sample_req_2061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(29), ack => phi_stmt_894_req_0); -- 
    -- Element group loadKernelChannel_CP_1909_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_entry_trigger
      -- 
    loadKernelChannel_CP_1909_elements(30) <= loadKernelChannel_CP_1909_elements(17);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_entry_sample_req_ps
      -- CP-element group 31: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_entry_sample_req
      -- 
    phi_stmt_894_entry_sample_req_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_894_entry_sample_req_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(31), ack => phi_stmt_894_req_1); -- 
    -- Element group loadKernelChannel_CP_1909_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_phi_mux_ack
      -- CP-element group 32: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_894_phi_mux_ack_ps
      -- 
    phi_stmt_894_phi_mux_ack_2067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_894_ack_0, ack => loadKernelChannel_CP_1909_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_Sample/req
      -- 
    req_2080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(33), ack => nmycount_916_896_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1909_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_Update/req
      -- CP-element group 34: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_update_start_
      -- CP-element group 34: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_update_start__ps
      -- 
    req_2085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(34), ack => nmycount_916_896_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1909_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_Sample/ack
      -- CP-element group 35: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_sample_completed__ps
      -- 
    ack_2081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_916_896_buf_ack_0, ack => loadKernelChannel_CP_1909_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nmycount_896_Update/$exit
      -- 
    ack_2086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_916_896_buf_ack_1, ack => loadKernelChannel_CP_1909_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_sample_start__ps
      -- 
    req_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(37), ack => start_add_897_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1909_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_update_start_
      -- CP-element group 38: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_Update/req
      -- 
    req_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(38), ack => start_add_897_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1909_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_sample_completed_
      -- 
    ack_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_897_buf_ack_0, ack => loadKernelChannel_CP_1909_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_start_add_897_Update/ack
      -- 
    ack_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_897_buf_ack_1, ack => loadKernelChannel_CP_1909_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	83 
    -- CP-element group 41: 	87 
    -- CP-element group 41: 	91 
    -- CP-element group 41: 	21 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_sample_start_
      -- 
    loadKernelChannel_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(18) & loadKernelChannel_CP_1909_elements(83) & loadKernelChannel_CP_1909_elements(87) & loadKernelChannel_CP_1909_elements(91) & loadKernelChannel_CP_1909_elements(21);
      gj_loadKernelChannel_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	64 
    -- CP-element group 42: 	67 
    -- CP-element group 42: 	90 
    -- CP-element group 42: 	46 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	22 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_update_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(18) & loadKernelChannel_CP_1909_elements(61) & loadKernelChannel_CP_1909_elements(64) & loadKernelChannel_CP_1909_elements(67) & loadKernelChannel_CP_1909_elements(90) & loadKernelChannel_CP_1909_elements(46);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_sample_start__ps
      -- 
    loadKernelChannel_CP_1909_elements(43) <= loadKernelChannel_CP_1909_elements(20);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1909_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_update_start__ps
      -- 
    loadKernelChannel_CP_1909_elements(45) <= loadKernelChannel_CP_1909_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	63 
    -- CP-element group 46: 	66 
    -- CP-element group 46: 	88 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_update_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1909_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_loopback_trigger
      -- 
    loadKernelChannel_CP_1909_elements(47) <= loadKernelChannel_CP_1909_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_loopback_sample_req
      -- CP-element group 48: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_loopback_sample_req_ps
      -- 
    phi_stmt_898_loopback_sample_req_2115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_898_loopback_sample_req_2115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(48), ack => phi_stmt_898_req_1); -- 
    -- Element group loadKernelChannel_CP_1909_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_entry_trigger
      -- 
    loadKernelChannel_CP_1909_elements(49) <= loadKernelChannel_CP_1909_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_entry_sample_req_ps
      -- 
    phi_stmt_898_entry_sample_req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_898_entry_sample_req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(50), ack => phi_stmt_898_req_0); -- 
    -- Element group loadKernelChannel_CP_1909_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/phi_stmt_898_phi_mux_ack_ps
      -- 
    phi_stmt_898_phi_mux_ack_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_898_ack_0, ack => loadKernelChannel_CP_1909_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_Sample/req
      -- 
    req_2134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(52), ack => my_fetch_861_900_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1909_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_update_start_
      -- CP-element group 53: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_Update/req
      -- 
    req_2139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(53), ack => my_fetch_861_900_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1909_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_Sample/ack
      -- 
    ack_2135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_861_900_buf_ack_0, ack => loadKernelChannel_CP_1909_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_my_fetch_900_Update/ack
      -- 
    ack_2140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_861_900_buf_ack_1, ack => loadKernelChannel_CP_1909_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_Sample/req
      -- 
    req_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(56), ack => nfetch_val_988_901_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1909_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_update_start_
      -- CP-element group 57: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_Update/req
      -- 
    req_2157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(57), ack => nfetch_val_988_901_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1909_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_sample_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_Sample/ack
      -- 
    ack_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_988_901_buf_ack_0, ack => loadKernelChannel_CP_1909_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_update_completed__ps
      -- CP-element group 59: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/R_nfetch_val_901_Update/ack
      -- 
    ack_2158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_988_901_buf_ack_1, ack => loadKernelChannel_CP_1909_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_Sample/req
      -- 
    req_2167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(60), ack => WPIPE_kernel_pipe1_942_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(27) & loadKernelChannel_CP_1909_elements(46) & loadKernelChannel_CP_1909_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	25 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_update_start_
      -- CP-element group 61: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_Update/req
      -- 
    ack_2168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_942_inst_ack_0, ack => loadKernelChannel_CP_1909_elements(61)); -- 
    req_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(61), ack => WPIPE_kernel_pipe1_942_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	93 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe1_942_Update/ack
      -- 
    ack_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_942_inst_ack_1, ack => loadKernelChannel_CP_1909_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	27 
    -- CP-element group 63: 	46 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_Sample/req
      -- 
    req_2181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(63), ack => WPIPE_kernel_pipe2_946_inst_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(27) & loadKernelChannel_CP_1909_elements(46) & loadKernelChannel_CP_1909_elements(65);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	25 
    -- CP-element group 64: 	42 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_update_start_
      -- CP-element group 64: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_Update/req
      -- 
    ack_2182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_946_inst_ack_0, ack => loadKernelChannel_CP_1909_elements(64)); -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(64), ack => WPIPE_kernel_pipe2_946_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	93 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe2_946_Update/ack
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_946_inst_ack_1, ack => loadKernelChannel_CP_1909_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	27 
    -- CP-element group 66: 	46 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_Sample/req
      -- 
    req_2195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(66), ack => WPIPE_kernel_pipe3_950_inst_req_0); -- 
    loadKernelChannel_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(27) & loadKernelChannel_CP_1909_elements(46) & loadKernelChannel_CP_1909_elements(68);
      gj_loadKernelChannel_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	42 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_update_start_
      -- CP-element group 67: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_Update/req
      -- 
    ack_2196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_950_inst_ack_0, ack => loadKernelChannel_CP_1909_elements(67)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(67), ack => WPIPE_kernel_pipe3_950_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	93 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/WPIPE_kernel_pipe3_950_Update/ack
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_950_inst_ack_1, ack => loadKernelChannel_CP_1909_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	73 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_request/$entry
      -- CP-element group 69: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_request/req
      -- 
    req_2241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(69), ack => addr_of_967_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(73) & loadKernelChannel_CP_1909_elements(74);
      gj_loadKernelChannel_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	18 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	75 
    -- CP-element group 70: 	82 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	75 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_update_start_
      -- CP-element group 70: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_complete/$entry
      -- CP-element group 70: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_complete/req
      -- 
    req_2246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(70), ack => addr_of_967_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(18) & loadKernelChannel_CP_1909_elements(75) & loadKernelChannel_CP_1909_elements(82);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	18 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	74 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_update_start
      -- CP-element group 71: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_Update/req
      -- 
    req_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(71), ack => array_obj_ref_966_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(18) & loadKernelChannel_CP_1909_elements(73) & loadKernelChannel_CP_1909_elements(74);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	27 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	93 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_sample_complete
      -- CP-element group 72: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_Sample/ack
      -- 
    ack_2227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_966_index_offset_ack_0, ack => loadKernelChannel_CP_1909_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (8) 
      -- CP-element group 73: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_offset_calculated
      -- CP-element group 73: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_final_index_sum_regn_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/array_obj_ref_966_base_plus_offset/sum_rename_ack
      -- 
    ack_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_966_index_offset_ack_1, ack => loadKernelChannel_CP_1909_elements(73)); -- 
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	71 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_request/$exit
      -- CP-element group 74: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_request/ack
      -- 
    ack_2242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_967_final_reg_ack_0, ack => loadKernelChannel_CP_1909_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	70 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	80 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	70 
    -- CP-element group 75:  members (19) 
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_word_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/addr_of_967_complete/ack
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_root_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_address_resized
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_addr_resize/$entry
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_addr_resize/$exit
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_addr_resize/base_resize_req
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_addr_resize/base_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_plus_offset/$entry
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_plus_offset/$exit
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_plus_offset/sum_rename_req
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_base_plus_offset/sum_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_word_addrgen/$entry
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_word_addrgen/$exit
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_word_addrgen/root_register_req
      -- CP-element group 75: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_word_addrgen/root_register_ack
      -- 
    ack_2247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_967_final_reg_ack_1, ack => loadKernelChannel_CP_1909_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	27 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_Sample/req
      -- 
    req_2255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(76), ack => W_fn_921_delayed_7_0_969_inst_req_0); -- 
    loadKernelChannel_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(27) & loadKernelChannel_CP_1909_elements(78);
      gj_loadKernelChannel_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	82 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_update_start_
      -- CP-element group 77: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_Update/req
      -- 
    req_2260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(77), ack => W_fn_921_delayed_7_0_969_inst_req_1); -- 
    loadKernelChannel_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(79) & loadKernelChannel_CP_1909_elements(82);
      gj_loadKernelChannel_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	25 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_Sample/ack
      -- 
    ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_921_delayed_7_0_969_inst_ack_0, ack => loadKernelChannel_CP_1909_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_971_Update/ack
      -- 
    ack_2261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_921_delayed_7_0_969_inst_ack_1, ack => loadKernelChannel_CP_1909_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: 	79 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Sample/word_access_start/word_0/rr
      -- 
    rr_2294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(80), ack => ptr_deref_975_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(75) & loadKernelChannel_CP_1909_elements(79) & loadKernelChannel_CP_1909_elements(82);
      gj_loadKernelChannel_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	21 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_update_start_
      -- CP-element group 81: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/word_access_complete/word_0/cr
      -- 
    cr_2305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(81), ack => ptr_deref_975_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(21) & loadKernelChannel_CP_1909_elements(83);
      gj_loadKernelChannel_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Sample/word_access_start/$exit
      -- CP-element group 82: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Sample/word_access_start/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Sample/word_access_start/word_0/ra
      -- 
    ra_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_975_load_0_ack_0, ack => loadKernelChannel_CP_1909_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	93 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	41 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/word_access_complete/$exit
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/word_access_complete/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/word_access_complete/word_0/ca
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/ptr_deref_975_Merge/$entry
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/ptr_deref_975_Merge/$exit
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/ptr_deref_975_Merge/merge_req
      -- CP-element group 83: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/ptr_deref_975_Update/ptr_deref_975_Merge/merge_ack
      -- 
    ca_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_975_load_0_ack_1, ack => loadKernelChannel_CP_1909_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	27 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_Sample/req
      -- 
    req_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(84), ack => W_fn_927_delayed_13_0_977_inst_req_0); -- 
    loadKernelChannel_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(27) & loadKernelChannel_CP_1909_elements(86);
      gj_loadKernelChannel_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	21 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_update_start_
      -- CP-element group 85: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_Update/req
      -- 
    req_2324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(85), ack => W_fn_927_delayed_13_0_977_inst_req_1); -- 
    loadKernelChannel_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(21) & loadKernelChannel_CP_1909_elements(87);
      gj_loadKernelChannel_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	25 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_Sample/ack
      -- 
    ack_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_927_delayed_13_0_977_inst_ack_0, ack => loadKernelChannel_CP_1909_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	93 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	41 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_979_Update/ack
      -- 
    ack_2325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_927_delayed_13_0_977_inst_ack_1, ack => loadKernelChannel_CP_1909_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	46 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_Sample/req
      -- 
    req_2333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(88), ack => W_fetch_val_929_delayed_13_0_980_inst_req_0); -- 
    loadKernelChannel_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(46) & loadKernelChannel_CP_1909_elements(90);
      gj_loadKernelChannel_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	21 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_update_start_
      -- CP-element group 89: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_Update/req
      -- 
    req_2338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(89), ack => W_fetch_val_929_delayed_13_0_980_inst_req_1); -- 
    loadKernelChannel_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(21) & loadKernelChannel_CP_1909_elements(91);
      gj_loadKernelChannel_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	42 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_Sample/ack
      -- 
    ack_2334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_929_delayed_13_0_980_inst_ack_0, ack => loadKernelChannel_CP_1909_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	41 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/assign_stmt_982_Update/ack
      -- 
    ack_2339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_929_delayed_13_0_980_inst_ack_1, ack => loadKernelChannel_CP_1909_elements(91)); -- 
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	18 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	19 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_1909_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_1909_elements(18), ack => loadKernelChannel_CP_1909_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	62 
    -- CP-element group 93: 	65 
    -- CP-element group 93: 	68 
    -- CP-element group 93: 	72 
    -- CP-element group 93: 	83 
    -- CP-element group 93: 	87 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	21 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	15 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_891/do_while_stmt_892/do_while_stmt_892_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1909_elements(62) & loadKernelChannel_CP_1909_elements(65) & loadKernelChannel_CP_1909_elements(68) & loadKernelChannel_CP_1909_elements(72) & loadKernelChannel_CP_1909_elements(83) & loadKernelChannel_CP_1909_elements(87) & loadKernelChannel_CP_1909_elements(91) & loadKernelChannel_CP_1909_elements(21);
      gj_loadKernelChannel_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_891/do_while_stmt_892/loop_exit/$exit
      -- CP-element group 94: 	 branch_block_stmt_891/do_while_stmt_892/loop_exit/ack
      -- 
    ack_2344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_892_branch_ack_0, ack => loadKernelChannel_CP_1909_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	14 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_891/do_while_stmt_892/loop_taken/$exit
      -- CP-element group 95: 	 branch_block_stmt_891/do_while_stmt_892/loop_taken/ack
      -- 
    ack_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_892_branch_ack_1, ack => loadKernelChannel_CP_1909_elements(95)); -- 
    -- CP-element group 96:  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	12 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	10 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_891/do_while_stmt_892/$exit
      -- 
    loadKernelChannel_CP_1909_elements(96) <= loadKernelChannel_CP_1909_elements(12);
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	10 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 assign_stmt_998/WPIPE_size_pipe_996_sample_completed_
      -- CP-element group 97: 	 assign_stmt_998/WPIPE_size_pipe_996_update_start_
      -- CP-element group 97: 	 assign_stmt_998/WPIPE_size_pipe_996_Sample/$exit
      -- CP-element group 97: 	 assign_stmt_998/WPIPE_size_pipe_996_Sample/ack
      -- CP-element group 97: 	 assign_stmt_998/WPIPE_size_pipe_996_Update/$entry
      -- CP-element group 97: 	 assign_stmt_998/WPIPE_size_pipe_996_Update/req
      -- 
    ack_2361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_996_inst_ack_0, ack => loadKernelChannel_CP_1909_elements(97)); -- 
    req_2365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1909_elements(97), ack => WPIPE_size_pipe_996_inst_req_1); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 $exit
      -- CP-element group 98: 	 assign_stmt_998/$exit
      -- CP-element group 98: 	 assign_stmt_998/WPIPE_size_pipe_996_update_completed_
      -- CP-element group 98: 	 assign_stmt_998/WPIPE_size_pipe_996_Update/$exit
      -- CP-element group 98: 	 assign_stmt_998/WPIPE_size_pipe_996_Update/ack
      -- 
    ack_2366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_996_inst_ack_1, ack => loadKernelChannel_CP_1909_elements(98)); -- 
    loadKernelChannel_do_while_stmt_892_terminator_2349: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_892_terminator_2349", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_1909_elements(15),loop_continue => loadKernelChannel_CP_1909_elements(95),loop_terminate => loadKernelChannel_CP_1909_elements(94),loop_back => loadKernelChannel_CP_1909_elements(13),loop_exit => loadKernelChannel_CP_1909_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_894_phi_seq_2105_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1909_elements(28);
      loadKernelChannel_CP_1909_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1909_elements(35);
      loadKernelChannel_CP_1909_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1909_elements(36);
      loadKernelChannel_CP_1909_elements(29) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1909_elements(30);
      loadKernelChannel_CP_1909_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1909_elements(39);
      loadKernelChannel_CP_1909_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1909_elements(40);
      loadKernelChannel_CP_1909_elements(31) <= phi_mux_reqs(1);
      phi_stmt_894_phi_seq_2105 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_894_phi_seq_2105") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1909_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_1909_elements(26), 
          phi_update_req => loadKernelChannel_CP_1909_elements(22), 
          phi_update_ack => loadKernelChannel_CP_1909_elements(27), 
          phi_mux_ack => loadKernelChannel_CP_1909_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_898_phi_seq_2159_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1909_elements(49);
      loadKernelChannel_CP_1909_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1909_elements(54);
      loadKernelChannel_CP_1909_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1909_elements(55);
      loadKernelChannel_CP_1909_elements(50) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1909_elements(47);
      loadKernelChannel_CP_1909_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1909_elements(58);
      loadKernelChannel_CP_1909_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1909_elements(59);
      loadKernelChannel_CP_1909_elements(48) <= phi_mux_reqs(1);
      phi_stmt_898_phi_seq_2159 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_898_phi_seq_2159") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1909_elements(43), 
          phi_sample_ack => loadKernelChannel_CP_1909_elements(44), 
          phi_update_req => loadKernelChannel_CP_1909_elements(45), 
          phi_update_ack => loadKernelChannel_CP_1909_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_1909_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2047_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_1909_elements(16);
        preds(1)  <= loadKernelChannel_CP_1909_elements(17);
        entry_tmerge_2047 : transition_merge -- 
          generic map(name => " entry_tmerge_2047")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_1909_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_907_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_956_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_920_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_965_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_965_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_965_wire : std_logic_vector(63 downto 0);
    signal NOT_u1_u1_930_wire : std_logic_vector(0 downto 0);
    signal R_sh_start_854_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_854_scaled : std_logic_vector(13 downto 0);
    signal SHL_u16_u16_843_wire : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_872_wire : std_logic_vector(15 downto 0);
    signal SUB_u64_u64_908_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_993_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_933_wire : std_logic_vector(0 downto 0);
    signal ULT_u64_u1_994_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_855_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_855_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_855_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_855_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_855_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_855_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_966_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_966_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_966_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_966_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_966_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_966_root_address : std_logic_vector(13 downto 0);
    signal ea1_867 : std_logic_vector(63 downto 0);
    signal ea2_875 : std_logic_vector(63 downto 0);
    signal ea3_881 : std_logic_vector(63 downto 0);
    signal fetch_addr_857 : std_logic_vector(31 downto 0);
    signal fetch_addr_968 : std_logic_vector(31 downto 0);
    signal fetch_val_898 : std_logic_vector(63 downto 0);
    signal fetch_val_929_delayed_13_0_982 : std_logic_vector(63 downto 0);
    signal first_fill_886 : std_logic_vector(0 downto 0);
    signal fn_921_delayed_7_0_971 : std_logic_vector(0 downto 0);
    signal fn_927_delayed_13_0_979 : std_logic_vector(0 downto 0);
    signal fn_959 : std_logic_vector(0 downto 0);
    signal fv_976 : std_logic_vector(63 downto 0);
    signal konst_842_wire_constant : std_logic_vector(15 downto 0);
    signal konst_848_wire_constant : std_logic_vector(63 downto 0);
    signal konst_871_wire_constant : std_logic_vector(15 downto 0);
    signal konst_884_wire_constant : std_logic_vector(63 downto 0);
    signal konst_904_wire_constant : std_logic_vector(63 downto 0);
    signal konst_906_wire_constant : std_logic_vector(63 downto 0);
    signal konst_909_wire_constant : std_logic_vector(63 downto 0);
    signal konst_914_wire_constant : std_logic_vector(63 downto 0);
    signal konst_955_wire_constant : std_logic_vector(63 downto 0);
    signal konst_957_wire_constant : std_logic_vector(63 downto 0);
    signal konst_964_wire_constant : std_logic_vector(63 downto 0);
    signal konst_992_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_861 : std_logic_vector(63 downto 0);
    signal my_fetch_861_900_buffered : std_logic_vector(63 downto 0);
    signal my_num1_911 : std_logic_vector(63 downto 0);
    signal mycount_894 : std_logic_vector(63 downto 0);
    signal nfetch_val_988 : std_logic_vector(63 downto 0);
    signal nfetch_val_988_901_buffered : std_logic_vector(63 downto 0);
    signal nmycount_916 : std_logic_vector(63 downto 0);
    signal nmycount_916_896_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_860_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_860_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_860_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_860_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_860_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_975_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_975_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_975_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_975_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_975_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_size_845 : std_logic_vector(15 downto 0);
    signal send_to_1_927 : std_logic_vector(0 downto 0);
    signal send_to_2_935 : std_logic_vector(0 downto 0);
    signal send_to_3_940 : std_logic_vector(0 downto 0);
    signal sh_start_850 : std_logic_vector(63 downto 0);
    signal start_add_897_buffered : std_logic_vector(63 downto 0);
    signal start_next_890 : std_logic_vector(7 downto 0);
    signal type_cast_865_wire : std_logic_vector(63 downto 0);
    signal type_cast_873_wire : std_logic_vector(63 downto 0);
    signal type_cast_879_wire : std_logic_vector(63 downto 0);
    signal var_val_922 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_855_constant_part_of_offset <= "00000000000000";
    array_obj_ref_855_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_855_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_855_resized_base_address <= "00000000000000";
    array_obj_ref_966_constant_part_of_offset <= "00000000000000";
    array_obj_ref_966_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_966_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_966_resized_base_address <= "00000000000000";
    konst_842_wire_constant <= "0000000000000001";
    konst_848_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_871_wire_constant <= "0000000000000001";
    konst_884_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_904_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_906_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_909_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_914_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_955_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_957_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_964_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_992_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_860_word_offset_0 <= "00000000000000";
    ptr_deref_975_word_offset_0 <= "00000000000000";
    phi_stmt_894: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_916_896_buffered & start_add_897_buffered;
      req <= phi_stmt_894_req_0 & phi_stmt_894_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_894",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_894_ack_0,
          idata => idata,
          odata => mycount_894,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_894
    phi_stmt_898: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch_861_900_buffered & nfetch_val_988_901_buffered;
      req <= phi_stmt_898_req_0 & phi_stmt_898_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_898",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_898_ack_0,
          idata => idata,
          odata => fetch_val_898,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_898
    -- flow-through select operator MUX_987_inst
    nfetch_val_988 <= fv_976 when (fn_927_delayed_13_0_979(0) /=  '0') else fetch_val_929_delayed_13_0_982;
    W_fetch_val_929_delayed_13_0_980_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_929_delayed_13_0_980_inst_req_0;
      W_fetch_val_929_delayed_13_0_980_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_929_delayed_13_0_980_inst_req_1;
      W_fetch_val_929_delayed_13_0_980_inst_ack_1<= rack(0);
      W_fetch_val_929_delayed_13_0_980_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_929_delayed_13_0_980_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_929_delayed_13_0_982,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_921_delayed_7_0_969_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_921_delayed_7_0_969_inst_req_0;
      W_fn_921_delayed_7_0_969_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_921_delayed_7_0_969_inst_req_1;
      W_fn_921_delayed_7_0_969_inst_ack_1<= rack(0);
      W_fn_921_delayed_7_0_969_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_921_delayed_7_0_969_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_959,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_921_delayed_7_0_971,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_927_delayed_13_0_977_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_927_delayed_13_0_977_inst_req_0;
      W_fn_927_delayed_13_0_977_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_927_delayed_13_0_977_inst_req_1;
      W_fn_927_delayed_13_0_977_inst_ack_1<= rack(0);
      W_fn_927_delayed_13_0_977_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_927_delayed_13_0_977_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_959,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_927_delayed_13_0_979,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_856_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_856_final_reg_req_0;
      addr_of_856_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_856_final_reg_req_1;
      addr_of_856_final_reg_ack_1<= rack(0);
      addr_of_856_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_856_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_855_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_857,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_967_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_967_final_reg_req_0;
      addr_of_967_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_967_final_reg_req_1;
      addr_of_967_final_reg_ack_1<= rack(0);
      addr_of_967_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_967_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_966_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_861_900_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_861_900_buf_req_0;
      my_fetch_861_900_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_861_900_buf_req_1;
      my_fetch_861_900_buf_ack_1<= rack(0);
      my_fetch_861_900_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_861_900_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_861_900_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_988_901_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_988_901_buf_req_0;
      nfetch_val_988_901_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_988_901_buf_req_1;
      nfetch_val_988_901_buf_ack_1<= rack(0);
      nfetch_val_988_901_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_988_901_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_988,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_988_901_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_916_896_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_916_896_buf_req_0;
      nmycount_916_896_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_916_896_buf_req_1;
      nmycount_916_896_buf_ack_1<= rack(0);
      nmycount_916_896_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_916_896_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_916,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_916_896_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_897_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_897_buf_req_0;
      start_add_897_buf_ack_0<= wack(0);
      rreq(0) <= start_add_897_buf_req_1;
      start_add_897_buf_ack_1<= rack(0);
      start_add_897_buf : InterlockBuffer generic map ( -- 
        name => "start_add_897_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_897_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_865_inst
    process(row_size_845) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_845(15 downto 0);
      type_cast_865_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_873_inst
    process(SHL_u16_u16_872_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := SHL_u16_u16_872_wire(15 downto 0);
      type_cast_873_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_879_inst
    process(row_size_845) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_845(15 downto 0);
      type_cast_879_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_921_inst
    process(LSHR_u64_u64_920_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_920_wire(15 downto 0);
      var_val_922 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_855_index_1_rename
    process(R_sh_start_854_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_854_resized;
      ov(13 downto 0) := iv;
      R_sh_start_854_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_855_index_1_resize
    process(sh_start_850) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_850;
      ov := iv(13 downto 0);
      R_sh_start_854_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_855_root_address_inst
    process(array_obj_ref_855_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_855_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_855_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_966_index_1_rename
    process(LSHR_u64_u64_965_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_965_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_965_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_966_index_1_resize
    process(LSHR_u64_u64_965_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_965_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_965_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_966_root_address_inst
    process(array_obj_ref_966_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_966_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_966_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_860_addr_0
    process(ptr_deref_860_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_860_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_860_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_860_base_resize
    process(fetch_addr_857) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_857;
      ov := iv(13 downto 0);
      ptr_deref_860_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_860_gather_scatter
    process(ptr_deref_860_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_860_data_0;
      ov(63 downto 0) := iv;
      my_fetch_861 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_860_root_address_inst
    process(ptr_deref_860_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_860_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_860_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_975_addr_0
    process(ptr_deref_975_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_975_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_975_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_975_base_resize
    process(fetch_addr_968) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_968;
      ov := iv(13 downto 0);
      ptr_deref_975_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_975_gather_scatter
    process(ptr_deref_975_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_975_data_0;
      ov(63 downto 0) := iv;
      fv_976 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_975_root_address_inst
    process(ptr_deref_975_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_975_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_975_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_892_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_994_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_892_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_892_branch_req_0,
          ack0 => do_while_stmt_892_branch_ack_0,
          ack1 => do_while_stmt_892_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_844_inst
    process(num_chl_buffer, SHL_u16_u16_843_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_chl_buffer, SHL_u16_u16_843_wire, tmp_var);
      row_size_845 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_866_inst
    process(start_add_buffer, type_cast_865_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_865_wire, tmp_var);
      ea1_867 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_874_inst
    process(start_add_buffer, type_cast_873_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_873_wire, tmp_var);
      ea2_875 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_880_inst
    process(ea2_875, type_cast_879_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ea2_875, type_cast_879_wire, tmp_var);
      ea3_881 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_915_inst
    process(mycount_894) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_894, konst_914_wire_constant, tmp_var);
      nmycount_916 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_934_inst
    process(NOT_u1_u1_930_wire, ULT_u64_u1_933_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_930_wire, ULT_u64_u1_933_wire, tmp_var);
      send_to_2_935 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_907_inst
    process(mycount_894) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_894, konst_906_wire_constant, tmp_var);
      AND_u64_u64_907_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_956_inst
    process(nmycount_916) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_916, konst_955_wire_constant, tmp_var);
      AND_u64_u64_956_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_885_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_884_wire_constant, tmp_var);
      first_fill_886 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_958_inst
    process(AND_u64_u64_956_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_956_wire, konst_957_wire_constant, tmp_var);
      fn_959 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_849_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_848_wire_constant, tmp_var);
      sh_start_850 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_920_inst
    process(fetch_val_898, my_num1_911) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_898, my_num1_911, tmp_var);
      LSHR_u64_u64_920_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_965_inst
    process(nmycount_916) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_916, konst_964_wire_constant, tmp_var);
      LSHR_u64_u64_965_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_930_inst
    process(send_to_1_927) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", send_to_1_927, tmp_var);
      NOT_u1_u1_930_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u16_u16_843_inst
    process(num_chl_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(num_chl_buffer, konst_842_wire_constant, tmp_var);
      SHL_u16_u16_843_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_872_inst
    process(row_size_845) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(row_size_845, konst_871_wire_constant, tmp_var);
      SHL_u16_u16_872_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_910_inst
    process(SUB_u64_u64_908_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_908_wire, konst_909_wire_constant, tmp_var);
      my_num1_911 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_908_inst
    process(konst_904_wire_constant, AND_u64_u64_907_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_904_wire_constant, AND_u64_u64_907_wire, tmp_var);
      SUB_u64_u64_908_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_993_inst
    process(ea3_881) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(ea3_881, konst_992_wire_constant, tmp_var);
      SUB_u64_u64_993_wire <= tmp_var; --
    end process;
    -- binary operator UGE_u64_u1_939_inst
    process(mycount_894, ea2_875) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(mycount_894, ea2_875, tmp_var);
      send_to_3_940 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_926_inst
    process(mycount_894, ea1_867) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_894, ea1_867, tmp_var);
      send_to_1_927 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_933_inst
    process(mycount_894, ea2_875) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_894, ea2_875, tmp_var);
      ULT_u64_u1_933_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_994_inst
    process(mycount_894, SUB_u64_u64_993_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_894, SUB_u64_u64_993_wire, tmp_var);
      ULT_u64_u1_994_wire <= tmp_var; --
    end process;
    -- shared split operator group (23) : array_obj_ref_855_index_offset 
    ApIntAdd_group_23: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_854_scaled;
      array_obj_ref_855_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_855_index_offset_req_0;
      array_obj_ref_855_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_855_index_offset_req_1;
      array_obj_ref_855_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_23_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : array_obj_ref_966_index_offset 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_965_scaled;
      array_obj_ref_966_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_966_index_offset_req_0;
      array_obj_ref_966_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_966_index_offset_req_1;
      array_obj_ref_966_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared load operator group (0) : ptr_deref_860_load_0 ptr_deref_975_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_860_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_975_load_0_req_0;
      ptr_deref_860_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_975_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_860_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_975_load_0_req_1;
      ptr_deref_860_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_975_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_921_delayed_7_0_971(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_860_word_address_0 & ptr_deref_975_word_address_0;
      ptr_deref_860_data_0 <= data_out(127 downto 64);
      ptr_deref_975_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_889_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_889_inst_req_0;
      RPIPE_input_done_pipe_889_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_889_inst_req_1;
      RPIPE_input_done_pipe_889_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_886(0);
      start_next_890 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_942_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_942_inst_req_0;
      WPIPE_kernel_pipe1_942_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_942_inst_req_1;
      WPIPE_kernel_pipe1_942_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_927(0);
      data_in <= var_val_922;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe2_946_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_946_inst_req_0;
      WPIPE_kernel_pipe2_946_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_946_inst_req_1;
      WPIPE_kernel_pipe2_946_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_935(0);
      data_in <= var_val_922;
      kernel_pipe2_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_kernel_pipe3_950_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe3_950_inst_req_0;
      WPIPE_kernel_pipe3_950_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe3_950_inst_req_1;
      WPIPE_kernel_pipe3_950_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_940(0);
      data_in <= var_val_922;
      kernel_pipe3_write_2_gI: SplitGuardInterface generic map(name => "kernel_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "kernel_pipe3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe3_pipe_write_req(0),
          oack => kernel_pipe3_pipe_write_ack(0),
          odata => kernel_pipe3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_size_pipe_996_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_996_inst_req_0;
      WPIPE_size_pipe_996_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_996_inst_req_1;
      WPIPE_size_pipe_996_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= num_chl_buffer;
      size_pipe_write_3_gI: SplitGuardInterface generic map(name => "size_pipe_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_3: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(63 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_2367_start: Boolean;
  signal sendB_CP_2367_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_1383_branch_ack_0 : boolean;
  signal addr_of_1062_final_reg_ack_0 : boolean;
  signal type_cast_1364_inst_req_1 : boolean;
  signal ptr_deref_1066_load_0_req_1 : boolean;
  signal addr_of_1062_final_reg_req_0 : boolean;
  signal type_cast_1364_inst_ack_1 : boolean;
  signal ptr_deref_1290_store_0_req_0 : boolean;
  signal type_cast_1080_inst_req_1 : boolean;
  signal type_cast_1080_inst_ack_1 : boolean;
  signal type_cast_1070_inst_ack_0 : boolean;
  signal type_cast_1080_inst_ack_0 : boolean;
  signal array_obj_ref_1441_final_reg_req_0 : boolean;
  signal ptr_deref_1374_store_0_req_1 : boolean;
  signal type_cast_1070_inst_req_0 : boolean;
  signal ptr_deref_1290_store_0_req_1 : boolean;
  signal type_cast_1364_inst_ack_0 : boolean;
  signal if_stmt_1015_branch_req_0 : boolean;
  signal addr_of_1062_final_reg_ack_1 : boolean;
  signal type_cast_1070_inst_req_1 : boolean;
  signal type_cast_1070_inst_ack_1 : boolean;
  signal ptr_deref_1290_store_0_ack_0 : boolean;
  signal if_stmt_1015_branch_ack_1 : boolean;
  signal type_cast_1364_inst_req_0 : boolean;
  signal if_stmt_1383_branch_ack_1 : boolean;
  signal ptr_deref_1353_store_0_req_1 : boolean;
  signal ptr_deref_1353_store_0_ack_1 : boolean;
  signal array_obj_ref_1441_final_reg_ack_1 : boolean;
  signal if_stmt_1015_branch_ack_0 : boolean;
  signal type_cast_1080_inst_req_0 : boolean;
  signal addr_of_1062_final_reg_req_1 : boolean;
  signal ptr_deref_1066_load_0_ack_0 : boolean;
  signal ptr_deref_1374_store_0_ack_1 : boolean;
  signal if_stmt_1383_branch_req_0 : boolean;
  signal array_obj_ref_1061_index_offset_ack_1 : boolean;
  signal array_obj_ref_1441_final_reg_req_1 : boolean;
  signal array_obj_ref_1061_index_offset_req_1 : boolean;
  signal array_obj_ref_1061_index_offset_ack_0 : boolean;
  signal array_obj_ref_1061_index_offset_req_0 : boolean;
  signal ptr_deref_1066_load_0_ack_1 : boolean;
  signal ptr_deref_1066_load_0_req_0 : boolean;
  signal array_obj_ref_1441_final_reg_ack_0 : boolean;
  signal type_cast_1322_inst_ack_1 : boolean;
  signal type_cast_1322_inst_req_1 : boolean;
  signal type_cast_1090_inst_req_0 : boolean;
  signal type_cast_1090_inst_ack_0 : boolean;
  signal type_cast_1090_inst_req_1 : boolean;
  signal type_cast_1090_inst_ack_1 : boolean;
  signal ptr_deref_1353_store_0_ack_0 : boolean;
  signal type_cast_1322_inst_ack_0 : boolean;
  signal type_cast_1322_inst_req_0 : boolean;
  signal type_cast_1100_inst_req_0 : boolean;
  signal type_cast_1343_inst_ack_1 : boolean;
  signal type_cast_1100_inst_ack_0 : boolean;
  signal type_cast_1100_inst_req_1 : boolean;
  signal type_cast_1343_inst_req_1 : boolean;
  signal type_cast_1100_inst_ack_1 : boolean;
  signal ptr_deref_1353_store_0_req_0 : boolean;
  signal type_cast_1110_inst_req_0 : boolean;
  signal type_cast_1110_inst_ack_0 : boolean;
  signal type_cast_1110_inst_req_1 : boolean;
  signal type_cast_1343_inst_ack_0 : boolean;
  signal type_cast_1110_inst_ack_1 : boolean;
  signal type_cast_1301_inst_ack_1 : boolean;
  signal type_cast_1301_inst_req_1 : boolean;
  signal type_cast_1343_inst_req_0 : boolean;
  signal type_cast_1120_inst_req_0 : boolean;
  signal type_cast_1120_inst_ack_0 : boolean;
  signal type_cast_1120_inst_req_1 : boolean;
  signal type_cast_1120_inst_ack_1 : boolean;
  signal ptr_deref_1311_store_0_ack_1 : boolean;
  signal ptr_deref_1311_store_0_req_1 : boolean;
  signal type_cast_1130_inst_req_0 : boolean;
  signal type_cast_1130_inst_ack_0 : boolean;
  signal type_cast_1130_inst_req_1 : boolean;
  signal type_cast_1130_inst_ack_1 : boolean;
  signal type_cast_1301_inst_ack_0 : boolean;
  signal type_cast_1140_inst_req_0 : boolean;
  signal type_cast_1140_inst_ack_0 : boolean;
  signal type_cast_1140_inst_req_1 : boolean;
  signal ptr_deref_1332_store_0_ack_1 : boolean;
  signal type_cast_1140_inst_ack_1 : boolean;
  signal type_cast_1301_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1142_inst_req_0 : boolean;
  signal ptr_deref_1332_store_0_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1142_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1142_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1142_inst_ack_1 : boolean;
  signal ptr_deref_1311_store_0_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1145_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1145_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1145_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1145_inst_ack_1 : boolean;
  signal ptr_deref_1311_store_0_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1148_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1148_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1148_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1148_inst_ack_1 : boolean;
  signal ptr_deref_1374_store_0_ack_0 : boolean;
  signal ptr_deref_1374_store_0_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1151_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1151_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1151_inst_req_1 : boolean;
  signal ptr_deref_1332_store_0_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1151_inst_ack_1 : boolean;
  signal array_obj_ref_1441_index_offset_ack_1 : boolean;
  signal array_obj_ref_1441_index_offset_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1154_inst_req_0 : boolean;
  signal ptr_deref_1332_store_0_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1154_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1154_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1154_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1157_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1157_inst_ack_0 : boolean;
  signal ptr_deref_1290_store_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1157_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1157_inst_ack_1 : boolean;
  signal array_obj_ref_1441_index_offset_ack_0 : boolean;
  signal array_obj_ref_1441_index_offset_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1160_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1160_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1160_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1160_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1163_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1163_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1163_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1163_inst_ack_1 : boolean;
  signal if_stmt_1177_branch_req_0 : boolean;
  signal if_stmt_1177_branch_ack_1 : boolean;
  signal if_stmt_1177_branch_ack_0 : boolean;
  signal if_stmt_1229_branch_req_0 : boolean;
  signal if_stmt_1229_branch_ack_1 : boolean;
  signal if_stmt_1229_branch_ack_0 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal array_obj_ref_1244_index_offset_req_0 : boolean;
  signal array_obj_ref_1244_index_offset_ack_0 : boolean;
  signal array_obj_ref_1244_index_offset_req_1 : boolean;
  signal array_obj_ref_1244_index_offset_ack_1 : boolean;
  signal addr_of_1245_final_reg_req_0 : boolean;
  signal addr_of_1245_final_reg_ack_0 : boolean;
  signal addr_of_1245_final_reg_req_1 : boolean;
  signal addr_of_1245_final_reg_ack_1 : boolean;
  signal ptr_deref_1249_load_0_req_0 : boolean;
  signal ptr_deref_1249_load_0_ack_0 : boolean;
  signal ptr_deref_1249_load_0_req_1 : boolean;
  signal ptr_deref_1249_load_0_ack_1 : boolean;
  signal type_cast_1259_inst_req_0 : boolean;
  signal type_cast_1259_inst_ack_0 : boolean;
  signal type_cast_1259_inst_req_1 : boolean;
  signal type_cast_1259_inst_ack_1 : boolean;
  signal ptr_deref_1269_store_0_req_0 : boolean;
  signal ptr_deref_1269_store_0_ack_0 : boolean;
  signal ptr_deref_1269_store_0_req_1 : boolean;
  signal ptr_deref_1269_store_0_ack_1 : boolean;
  signal type_cast_1280_inst_req_0 : boolean;
  signal type_cast_1280_inst_ack_0 : boolean;
  signal type_cast_1280_inst_req_1 : boolean;
  signal type_cast_1280_inst_ack_1 : boolean;
  signal array_obj_ref_1453_index_offset_req_0 : boolean;
  signal array_obj_ref_1453_index_offset_ack_0 : boolean;
  signal array_obj_ref_1453_index_offset_req_1 : boolean;
  signal array_obj_ref_1453_index_offset_ack_1 : boolean;
  signal array_obj_ref_1453_final_reg_req_0 : boolean;
  signal array_obj_ref_1453_final_reg_ack_0 : boolean;
  signal array_obj_ref_1453_final_reg_req_1 : boolean;
  signal array_obj_ref_1453_final_reg_ack_1 : boolean;
  signal ptr_deref_1457_load_0_req_0 : boolean;
  signal ptr_deref_1457_load_0_ack_0 : boolean;
  signal ptr_deref_1457_load_0_req_1 : boolean;
  signal ptr_deref_1457_load_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1459_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1459_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1459_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1459_inst_ack_1 : boolean;
  signal ptr_deref_1464_load_0_req_0 : boolean;
  signal ptr_deref_1464_load_0_ack_0 : boolean;
  signal ptr_deref_1464_load_0_req_1 : boolean;
  signal ptr_deref_1464_load_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1466_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1466_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1466_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1466_inst_ack_1 : boolean;
  signal if_stmt_1480_branch_req_0 : boolean;
  signal if_stmt_1480_branch_ack_1 : boolean;
  signal if_stmt_1480_branch_ack_0 : boolean;
  signal phi_stmt_1049_req_0 : boolean;
  signal type_cast_1055_inst_req_0 : boolean;
  signal type_cast_1055_inst_ack_0 : boolean;
  signal type_cast_1055_inst_req_1 : boolean;
  signal type_cast_1055_inst_ack_1 : boolean;
  signal phi_stmt_1049_req_1 : boolean;
  signal phi_stmt_1049_ack_0 : boolean;
  signal phi_stmt_1209_req_1 : boolean;
  signal type_cast_1212_inst_req_0 : boolean;
  signal type_cast_1212_inst_ack_0 : boolean;
  signal type_cast_1212_inst_req_1 : boolean;
  signal type_cast_1212_inst_ack_1 : boolean;
  signal phi_stmt_1209_req_0 : boolean;
  signal phi_stmt_1209_ack_0 : boolean;
  signal phi_stmt_1423_req_0 : boolean;
  signal type_cast_1429_inst_req_0 : boolean;
  signal type_cast_1429_inst_ack_0 : boolean;
  signal type_cast_1429_inst_req_1 : boolean;
  signal type_cast_1429_inst_ack_1 : boolean;
  signal phi_stmt_1423_req_1 : boolean;
  signal phi_stmt_1423_ack_0 : boolean;
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= size;
  size_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_2367_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2367_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_2367_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2367_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_2367: Block -- control-path 
    signal sendB_CP_2367_elements: BooleanArray(137 downto 0);
    -- 
  begin -- 
    sendB_CP_2367_elements(0) <= sendB_CP_2367_start;
    sendB_CP_2367_symbol <= sendB_CP_2367_elements(137);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_1002/if_stmt_1015__entry__
      -- CP-element group 0: 	 branch_block_stmt_1002/assign_stmt_1008_to_assign_stmt_1014/$entry
      -- CP-element group 0: 	 branch_block_stmt_1002/assign_stmt_1008_to_assign_stmt_1014__exit__
      -- CP-element group 0: 	 branch_block_stmt_1002/if_stmt_1015_else_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1002/assign_stmt_1008_to_assign_stmt_1014/$exit
      -- CP-element group 0: 	 branch_block_stmt_1002/if_stmt_1015_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1002/if_stmt_1015_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_1002/if_stmt_1015_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_1002/if_stmt_1015_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1002/if_stmt_1015_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_1002/assign_stmt_1008_to_assign_stmt_1014__entry__
      -- CP-element group 0: 	 branch_block_stmt_1002/R_cmp77_1016_place
      -- CP-element group 0: 	 branch_block_stmt_1002/branch_block_stmt_1002__entry__
      -- CP-element group 0: 	 branch_block_stmt_1002/$entry
      -- CP-element group 0: 	 $entry
      -- 
    branch_req_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(0), ack => if_stmt_1015_branch_req_0); -- 
    -- CP-element group 1:  merge  transition  place  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	119 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_1002/merge_stmt_1021__exit__
      -- CP-element group 1: 	 branch_block_stmt_1002/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_1002/assign_stmt_1027_to_assign_stmt_1046/$entry
      -- CP-element group 1: 	 branch_block_stmt_1002/if_stmt_1015_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody
      -- CP-element group 1: 	 branch_block_stmt_1002/assign_stmt_1027_to_assign_stmt_1046__exit__
      -- CP-element group 1: 	 branch_block_stmt_1002/assign_stmt_1027_to_assign_stmt_1046__entry__
      -- CP-element group 1: 	 branch_block_stmt_1002/if_stmt_1015_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_1002/assign_stmt_1027_to_assign_stmt_1046/$exit
      -- CP-element group 1: 	 branch_block_stmt_1002/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1002/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_1002/merge_stmt_1021_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_1002/merge_stmt_1021_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_1002/merge_stmt_1021_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_1002/merge_stmt_1021_PhiAck/dummy
      -- CP-element group 1: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1049/$entry
      -- CP-element group 1: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/$entry
      -- 
    if_choice_transition_2436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1015_branch_ack_1, ack => sendB_CP_2367_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	125 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1002/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_1002/if_stmt_1015_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_1002/if_stmt_1015_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_1002/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1002/entry_forx_xend_PhiReq/phi_stmt_1209/$entry
      -- CP-element group 2: 	 branch_block_stmt_1002/entry_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/$entry
      -- 
    else_choice_transition_2440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1015_branch_ack_0, ack => sendB_CP_2367_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	124 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	48 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_sample_complete
      -- CP-element group 3: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_Sample/ack
      -- 
    ack_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1061_index_offset_ack_0, ack => sendB_CP_2367_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	124 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (11) 
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_request/$entry
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_request/req
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_offset_calculated
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_base_plus_offset/$entry
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_base_plus_offset/$exit
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_root_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_Update/ack
      -- CP-element group 4: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_Update/$exit
      -- 
    ack_2479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1061_index_offset_ack_1, ack => sendB_CP_2367_elements(4)); -- 
    req_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(4), ack => addr_of_1062_final_reg_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_request/$exit
      -- CP-element group 5: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_request/ack
      -- CP-element group 5: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_sample_completed_
      -- 
    ack_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1062_final_reg_ack_0, ack => sendB_CP_2367_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	124 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (24) 
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_word_addrgen/$entry
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_word_addrgen/root_register_ack
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_addr_resize/base_resize_req
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_word_addrgen/$exit
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_complete/ack
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_addr_resize/base_resize_ack
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_address_resized
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_word_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_addr_resize/$exit
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_word_addrgen/root_register_req
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Sample/word_access_start/$entry
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Sample/word_access_start/word_0/rr
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_base_addr_resize/$entry
      -- CP-element group 6: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Sample/$entry
      -- 
    ack_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1062_final_reg_ack_1, ack => sendB_CP_2367_elements(6)); -- 
    rr_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(6), ack => ptr_deref_1066_load_0_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Sample/word_access_start/word_0/ra
      -- 
    ra_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1066_load_0_ack_0, ack => sendB_CP_2367_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	124 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	15 
    -- CP-element group 8: 	17 
    -- CP-element group 8: 	19 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	11 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (33) 
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/ptr_deref_1066_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/ptr_deref_1066_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/ptr_deref_1066_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/ptr_deref_1066_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_Sample/rr
      -- 
    ca_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1066_load_0_ack_1, ack => sendB_CP_2367_elements(8)); -- 
    rr_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(8), ack => type_cast_1070_inst_req_0); -- 
    rr_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(8), ack => type_cast_1110_inst_req_0); -- 
    rr_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(8), ack => type_cast_1120_inst_req_0); -- 
    rr_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(8), ack => type_cast_1130_inst_req_0); -- 
    rr_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(8), ack => type_cast_1140_inst_req_0); -- 
    rr_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(8), ack => type_cast_1080_inst_req_0); -- 
    rr_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(8), ack => type_cast_1090_inst_req_0); -- 
    rr_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(8), ack => type_cast_1100_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_sample_completed_
      -- 
    ra_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1070_inst_ack_0, ack => sendB_CP_2367_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	124 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	45 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_Update/ca
      -- 
    ca_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1070_inst_ack_1, ack => sendB_CP_2367_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_Sample/$exit
      -- 
    ra_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1080_inst_ack_0, ack => sendB_CP_2367_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	124 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	42 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_Update/$exit
      -- 
    ca_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1080_inst_ack_1, ack => sendB_CP_2367_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_Sample/ra
      -- 
    ra_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1090_inst_ack_0, ack => sendB_CP_2367_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	124 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	39 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_Update/ca
      -- 
    ca_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1090_inst_ack_1, ack => sendB_CP_2367_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	8 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_Sample/ra
      -- 
    ra_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1100_inst_ack_0, ack => sendB_CP_2367_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	124 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	36 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_Update/ca
      -- 
    ca_2600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1100_inst_ack_1, ack => sendB_CP_2367_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	8 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_Sample/ra
      -- 
    ra_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_0, ack => sendB_CP_2367_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	124 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_Update/ca
      -- 
    ca_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_1, ack => sendB_CP_2367_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	8 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_Sample/ra
      -- 
    ra_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1120_inst_ack_0, ack => sendB_CP_2367_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	124 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	30 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_Update/ca
      -- 
    ca_2628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1120_inst_ack_1, ack => sendB_CP_2367_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_Sample/ra
      -- 
    ra_2637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_0, ack => sendB_CP_2367_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	124 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_Update/ca
      -- 
    ca_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_1, ack => sendB_CP_2367_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_Sample/ra
      -- 
    ra_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1140_inst_ack_0, ack => sendB_CP_2367_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	124 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_Sample/req
      -- 
    ca_2656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1140_inst_ack_1, ack => sendB_CP_2367_elements(24)); -- 
    req_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(24), ack => WPIPE_maxpool_output_pipe_1142_inst_req_0); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_Sample/ack
      -- CP-element group 25: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_Update/req
      -- 
    ack_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1142_inst_ack_0, ack => sendB_CP_2367_elements(25)); -- 
    req_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(25), ack => WPIPE_maxpool_output_pipe_1142_inst_req_1); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1142_Update/ack
      -- 
    ack_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1142_inst_ack_1, ack => sendB_CP_2367_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: 	22 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_Sample/req
      -- 
    req_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(27), ack => WPIPE_maxpool_output_pipe_1145_inst_req_0); -- 
    sendB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(26) & sendB_CP_2367_elements(22);
      gj_sendB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_Update/req
      -- 
    ack_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1145_inst_ack_0, ack => sendB_CP_2367_elements(28)); -- 
    req_2683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(28), ack => WPIPE_maxpool_output_pipe_1145_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1145_Update/ack
      -- 
    ack_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1145_inst_ack_1, ack => sendB_CP_2367_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: 	20 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_Sample/req
      -- 
    req_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(30), ack => WPIPE_maxpool_output_pipe_1148_inst_req_0); -- 
    sendB_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(29) & sendB_CP_2367_elements(20);
      gj_sendB_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_Update/req
      -- 
    ack_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1148_inst_ack_0, ack => sendB_CP_2367_elements(31)); -- 
    req_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(31), ack => WPIPE_maxpool_output_pipe_1148_inst_req_1); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1148_Update/ack
      -- 
    ack_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1148_inst_ack_1, ack => sendB_CP_2367_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	18 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_Sample/req
      -- 
    req_2706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(33), ack => WPIPE_maxpool_output_pipe_1151_inst_req_0); -- 
    sendB_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(32) & sendB_CP_2367_elements(18);
      gj_sendB_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_Update/req
      -- 
    ack_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1151_inst_ack_0, ack => sendB_CP_2367_elements(34)); -- 
    req_2711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(34), ack => WPIPE_maxpool_output_pipe_1151_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1151_Update/ack
      -- 
    ack_2712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1151_inst_ack_1, ack => sendB_CP_2367_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	16 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_Sample/req
      -- 
    req_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(36), ack => WPIPE_maxpool_output_pipe_1154_inst_req_0); -- 
    sendB_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(35) & sendB_CP_2367_elements(16);
      gj_sendB_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_Update/req
      -- 
    ack_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1154_inst_ack_0, ack => sendB_CP_2367_elements(37)); -- 
    req_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(37), ack => WPIPE_maxpool_output_pipe_1154_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1154_Update/ack
      -- 
    ack_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1154_inst_ack_1, ack => sendB_CP_2367_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: 	14 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_Sample/req
      -- 
    req_2734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(39), ack => WPIPE_maxpool_output_pipe_1157_inst_req_0); -- 
    sendB_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(38) & sendB_CP_2367_elements(14);
      gj_sendB_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_Update/req
      -- 
    ack_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1157_inst_ack_0, ack => sendB_CP_2367_elements(40)); -- 
    req_2739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(40), ack => WPIPE_maxpool_output_pipe_1157_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1157_Update/ack
      -- 
    ack_2740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1157_inst_ack_1, ack => sendB_CP_2367_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	12 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_Sample/req
      -- 
    req_2748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(42), ack => WPIPE_maxpool_output_pipe_1160_inst_req_0); -- 
    sendB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(41) & sendB_CP_2367_elements(12);
      gj_sendB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_Update/req
      -- 
    ack_2749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1160_inst_ack_0, ack => sendB_CP_2367_elements(43)); -- 
    req_2753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(43), ack => WPIPE_maxpool_output_pipe_1160_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1160_Update/ack
      -- 
    ack_2754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1160_inst_ack_1, ack => sendB_CP_2367_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_Sample/req
      -- 
    req_2762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(45), ack => WPIPE_maxpool_output_pipe_1163_inst_req_0); -- 
    sendB_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(44) & sendB_CP_2367_elements(10);
      gj_sendB_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_Update/req
      -- 
    ack_2763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1163_inst_ack_0, ack => sendB_CP_2367_elements(46)); -- 
    req_2767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(46), ack => WPIPE_maxpool_output_pipe_1163_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/WPIPE_maxpool_output_pipe_1163_Update/ack
      -- 
    ack_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1163_inst_ack_1, ack => sendB_CP_2367_elements(47)); -- 
    -- CP-element group 48:  branch  join  transition  place  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	3 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (10) 
      -- CP-element group 48: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176__exit__
      -- CP-element group 48: 	 branch_block_stmt_1002/if_stmt_1177__entry__
      -- CP-element group 48: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/$exit
      -- CP-element group 48: 	 branch_block_stmt_1002/if_stmt_1177_dead_link/$entry
      -- CP-element group 48: 	 branch_block_stmt_1002/if_stmt_1177_eval_test/$entry
      -- CP-element group 48: 	 branch_block_stmt_1002/if_stmt_1177_eval_test/$exit
      -- CP-element group 48: 	 branch_block_stmt_1002/if_stmt_1177_eval_test/branch_req
      -- CP-element group 48: 	 branch_block_stmt_1002/R_exitcond_1178_place
      -- CP-element group 48: 	 branch_block_stmt_1002/if_stmt_1177_if_link/$entry
      -- CP-element group 48: 	 branch_block_stmt_1002/if_stmt_1177_else_link/$entry
      -- 
    branch_req_2776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(48), ack => if_stmt_1177_branch_req_0); -- 
    sendB_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(47) & sendB_CP_2367_elements(3);
      gj_sendB_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	126 
    -- CP-element group 49: 	127 
    -- CP-element group 49:  members (24) 
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 49: 	 branch_block_stmt_1002/assign_stmt_1190_to_assign_stmt_1206__exit__
      -- CP-element group 49: 	 branch_block_stmt_1002/assign_stmt_1190_to_assign_stmt_1206__entry__
      -- CP-element group 49: 	 branch_block_stmt_1002/merge_stmt_1183__exit__
      -- CP-element group 49: 	 branch_block_stmt_1002/if_stmt_1177_if_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_1002/if_stmt_1177_if_link/if_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 49: 	 branch_block_stmt_1002/assign_stmt_1190_to_assign_stmt_1206/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/assign_stmt_1190_to_assign_stmt_1206/$exit
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 49: 	 branch_block_stmt_1002/merge_stmt_1183_PhiReqMerge
      -- CP-element group 49: 	 branch_block_stmt_1002/merge_stmt_1183_PhiAck/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/merge_stmt_1183_PhiAck/$exit
      -- CP-element group 49: 	 branch_block_stmt_1002/merge_stmt_1183_PhiAck/dummy
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1177_branch_ack_1, ack => sendB_CP_2367_elements(49)); -- 
    rr_3676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(49), ack => type_cast_1212_inst_req_0); -- 
    cr_3681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(49), ack => type_cast_1212_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  place  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	120 
    -- CP-element group 50: 	121 
    -- CP-element group 50:  members (12) 
      -- CP-element group 50: 	 branch_block_stmt_1002/if_stmt_1177_else_link/$exit
      -- CP-element group 50: 	 branch_block_stmt_1002/if_stmt_1177_else_link/else_choice_transition
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/$entry
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/$entry
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/$entry
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/$entry
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1177_branch_ack_0, ack => sendB_CP_2367_elements(50)); -- 
    rr_3622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(50), ack => type_cast_1055_inst_req_0); -- 
    cr_3627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(50), ack => type_cast_1055_inst_req_1); -- 
    -- CP-element group 51:  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	130 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	137 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1002/if_stmt_1229_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_1002/if_stmt_1229_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_1002/forx_xend_sendRemainingElementsx_xexit
      -- CP-element group 51: 	 branch_block_stmt_1002/forx_xend_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1002/forx_xend_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_2806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1229_branch_ack_1, ack => sendB_CP_2367_elements(51)); -- 
    -- CP-element group 52:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	130 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	85 
    -- CP-element group 52: 	87 
    -- CP-element group 52: 	88 
    -- CP-element group 52: 	90 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52: 	56 
    -- CP-element group 52: 	58 
    -- CP-element group 52: 	75 
    -- CP-element group 52: 	77 
    -- CP-element group 52: 	78 
    -- CP-element group 52: 	80 
    -- CP-element group 52: 	82 
    -- CP-element group 52: 	83 
    -- CP-element group 52: 	67 
    -- CP-element group 52: 	68 
    -- CP-element group 52: 	70 
    -- CP-element group 52: 	72 
    -- CP-element group 52: 	73 
    -- CP-element group 52: 	60 
    -- CP-element group 52: 	62 
    -- CP-element group 52: 	63 
    -- CP-element group 52: 	65 
    -- CP-element group 52:  members (186) 
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/merge_stmt_1235__exit__
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382__entry__
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/if_stmt_1229_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/if_stmt_1229_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_1002/forx_xend_ifx_xthen
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_resized_1
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_scaled_1
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_computed_1
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_resize_1/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_resize_1/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_resize_1/index_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_resize_1/index_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_scale_1/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_scale_1/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_scale_1/scale_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_index_scale_1/scale_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_update_start
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_Update/req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_complete/req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1002/forx_xend_ifx_xthen_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/forx_xend_ifx_xthen_PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/merge_stmt_1235_PhiReqMerge
      -- CP-element group 52: 	 branch_block_stmt_1002/merge_stmt_1235_PhiAck/$entry
      -- CP-element group 52: 	 branch_block_stmt_1002/merge_stmt_1235_PhiAck/$exit
      -- CP-element group 52: 	 branch_block_stmt_1002/merge_stmt_1235_PhiAck/dummy
      -- 
    else_choice_transition_2810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1229_branch_ack_0, ack => sendB_CP_2367_elements(52)); -- 
    cr_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => type_cast_1364_inst_req_1); -- 
    cr_3308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => ptr_deref_1374_store_0_req_1); -- 
    cr_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => ptr_deref_1290_store_0_req_1); -- 
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => ptr_deref_1353_store_0_req_1); -- 
    cr_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => type_cast_1322_inst_req_1); -- 
    cr_3194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => type_cast_1343_inst_req_1); -- 
    cr_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => type_cast_1301_inst_req_1); -- 
    cr_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => ptr_deref_1311_store_0_req_1); -- 
    cr_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => ptr_deref_1332_store_0_req_1); -- 
    rr_2823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => type_cast_1238_inst_req_0); -- 
    cr_2828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => type_cast_1238_inst_req_1); -- 
    req_2854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => array_obj_ref_1244_index_offset_req_0); -- 
    req_2859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => array_obj_ref_1244_index_offset_req_1); -- 
    req_2874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => addr_of_1245_final_reg_req_1); -- 
    cr_2919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => ptr_deref_1249_load_0_req_1); -- 
    cr_2938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => type_cast_1259_inst_req_1); -- 
    cr_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => ptr_deref_1269_store_0_req_1); -- 
    cr_3002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(52), ack => type_cast_1280_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_Sample/ra
      -- 
    ra_2824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => sendB_CP_2367_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	96 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1238_Update/ca
      -- 
    ca_2829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => sendB_CP_2367_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	96 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_sample_complete
      -- CP-element group 55: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_Sample/ack
      -- 
    ack_2855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1244_index_offset_ack_0, ack => sendB_CP_2367_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	52 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (11) 
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_offset_calculated
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_final_index_sum_regn_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/array_obj_ref_1244_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_request/$entry
      -- CP-element group 56: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_request/req
      -- 
    ack_2860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1244_index_offset_ack_1, ack => sendB_CP_2367_elements(56)); -- 
    req_2869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(56), ack => addr_of_1245_final_reg_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_request/$exit
      -- CP-element group 57: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_request/ack
      -- 
    ack_2870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1245_final_reg_ack_0, ack => sendB_CP_2367_elements(57)); -- 
    -- CP-element group 58:  join  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	52 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_complete/$exit
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/addr_of_1245_complete/ack
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_address_resized
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_addr_resize/$entry
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_addr_resize/$exit
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_addr_resize/base_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_addr_resize/base_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_word_addrgen/$entry
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_word_addrgen/$exit
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_word_addrgen/root_register_req
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_word_addrgen/root_register_ack
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Sample/word_access_start/word_0/rr
      -- 
    ack_2875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1245_final_reg_ack_1, ack => sendB_CP_2367_elements(58)); -- 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(58), ack => ptr_deref_1249_load_0_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Sample/word_access_start/$exit
      -- CP-element group 59: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Sample/word_access_start/word_0/ra
      -- 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1249_load_0_ack_0, ack => sendB_CP_2367_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	52 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	86 
    -- CP-element group 60: 	76 
    -- CP-element group 60: 	81 
    -- CP-element group 60: 	66 
    -- CP-element group 60: 	71 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (27) 
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/word_access_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/ptr_deref_1249_Merge/$entry
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/ptr_deref_1249_Merge/$exit
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/ptr_deref_1249_Merge/merge_req
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1249_Update/ptr_deref_1249_Merge/merge_ack
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_Sample/rr
      -- 
    ca_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1249_load_0_ack_1, ack => sendB_CP_2367_elements(60)); -- 
    rr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(60), ack => type_cast_1364_inst_req_0); -- 
    rr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(60), ack => type_cast_1322_inst_req_0); -- 
    rr_3189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(60), ack => type_cast_1343_inst_req_0); -- 
    rr_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(60), ack => type_cast_1301_inst_req_0); -- 
    rr_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(60), ack => type_cast_1259_inst_req_0); -- 
    rr_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(60), ack => type_cast_1280_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_Sample/ra
      -- 
    ra_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_0, ack => sendB_CP_2367_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	52 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1259_Update/ca
      -- 
    ca_2939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_1, ack => sendB_CP_2367_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	52 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/ptr_deref_1269_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/ptr_deref_1269_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/ptr_deref_1269_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/ptr_deref_1269_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/word_access_start/word_0/rr
      -- 
    rr_2977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(63), ack => ptr_deref_1269_store_0_req_0); -- 
    sendB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(52) & sendB_CP_2367_elements(62);
      gj_sendB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	91 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Sample/word_access_start/word_0/ra
      -- 
    ra_2978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1269_store_0_ack_0, ack => sendB_CP_2367_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	52 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	96 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_Update/word_access_complete/word_0/ca
      -- 
    ca_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1269_store_0_ack_1, ack => sendB_CP_2367_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_Sample/ra
      -- 
    ra_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1280_inst_ack_0, ack => sendB_CP_2367_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	52 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1280_Update/ca
      -- 
    ca_3003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1280_inst_ack_1, ack => sendB_CP_2367_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	91 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (9) 
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/word_access_start/$entry
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/word_access_start/word_0/rr
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/word_access_start/word_0/$entry
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/ptr_deref_1290_Split/$entry
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/ptr_deref_1290_Split/split_ack
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/ptr_deref_1290_Split/split_req
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/ptr_deref_1290_Split/$exit
      -- CP-element group 68: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_sample_start_
      -- 
    rr_3041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(68), ack => ptr_deref_1290_store_0_req_0); -- 
    sendB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(91) & sendB_CP_2367_elements(52) & sendB_CP_2367_elements(67);
      gj_sendB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	92 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/word_access_start/$exit
      -- CP-element group 69: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/word_access_start/word_0/ra
      -- CP-element group 69: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Sample/word_access_start/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_sample_completed_
      -- 
    ra_3042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1290_store_0_ack_0, ack => sendB_CP_2367_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	52 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	96 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Update/word_access_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Update/word_access_complete/word_0/$exit
      -- CP-element group 70: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_Update/word_access_complete/word_0/ca
      -- 
    ca_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1290_store_0_ack_1, ack => sendB_CP_2367_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	60 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_sample_completed_
      -- 
    ra_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1301_inst_ack_0, ack => sendB_CP_2367_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	52 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1301_update_completed_
      -- 
    ca_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1301_inst_ack_1, ack => sendB_CP_2367_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	92 
    -- CP-element group 73: 	52 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/ptr_deref_1311_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/ptr_deref_1311_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/ptr_deref_1311_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/ptr_deref_1311_Split/split_ack
      -- 
    rr_3105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(73), ack => ptr_deref_1311_store_0_req_0); -- 
    sendB_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(92) & sendB_CP_2367_elements(52) & sendB_CP_2367_elements(72);
      gj_sendB_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	93 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/word_access_start/word_0/ra
      -- CP-element group 74: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Sample/word_access_start/$exit
      -- 
    ra_3106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1311_store_0_ack_0, ack => sendB_CP_2367_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	96 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Update/word_access_complete/word_0/ca
      -- CP-element group 75: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_Update/$exit
      -- 
    ca_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1311_store_0_ack_1, ack => sendB_CP_2367_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	60 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_sample_completed_
      -- 
    ra_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1322_inst_ack_0, ack => sendB_CP_2367_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	52 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1322_update_completed_
      -- 
    ca_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1322_inst_ack_1, ack => sendB_CP_2367_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	93 
    -- CP-element group 78: 	52 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/ptr_deref_1332_Split/$exit
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/ptr_deref_1332_Split/$entry
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/ptr_deref_1332_Split/split_req
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/ptr_deref_1332_Split/split_ack
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/word_access_start/$entry
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/word_access_start/word_0/rr
      -- CP-element group 78: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/word_access_start/word_0/$entry
      -- 
    rr_3169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(78), ack => ptr_deref_1332_store_0_req_0); -- 
    sendB_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(93) & sendB_CP_2367_elements(52) & sendB_CP_2367_elements(77);
      gj_sendB_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	94 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/word_access_start/word_0/ra
      -- CP-element group 79: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/word_access_start/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Sample/word_access_start/$exit
      -- 
    ra_3170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1332_store_0_ack_0, ack => sendB_CP_2367_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	52 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	96 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Update/word_access_complete/word_0/ca
      -- CP-element group 80: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Update/word_access_complete/word_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Update/word_access_complete/$exit
      -- CP-element group 80: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_Update/$exit
      -- 
    ca_3181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1332_store_0_ack_1, ack => sendB_CP_2367_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	60 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_sample_completed_
      -- 
    ra_3190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1343_inst_ack_0, ack => sendB_CP_2367_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	52 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1343_update_completed_
      -- 
    ca_3195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1343_inst_ack_1, ack => sendB_CP_2367_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	94 
    -- CP-element group 83: 	52 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/word_access_start/word_0/rr
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/word_access_start/word_0/$entry
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/word_access_start/$entry
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/ptr_deref_1353_Split/split_ack
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/ptr_deref_1353_Split/split_req
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/ptr_deref_1353_Split/$exit
      -- CP-element group 83: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/ptr_deref_1353_Split/$entry
      -- 
    rr_3233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(83), ack => ptr_deref_1353_store_0_req_0); -- 
    sendB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(94) & sendB_CP_2367_elements(52) & sendB_CP_2367_elements(82);
      gj_sendB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	95 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/word_access_start/word_0/ra
      -- CP-element group 84: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/word_access_start/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Sample/word_access_start/$exit
      -- 
    ra_3234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1353_store_0_ack_0, ack => sendB_CP_2367_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	52 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	96 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Update/word_access_complete/$exit
      -- CP-element group 85: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Update/word_access_complete/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Update/word_access_complete/word_0/ca
      -- CP-element group 85: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_Update/$exit
      -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1353_store_0_ack_1, ack => sendB_CP_2367_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	60 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_Sample/$exit
      -- 
    ra_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1364_inst_ack_0, ack => sendB_CP_2367_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	52 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/type_cast_1364_update_completed_
      -- 
    ca_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1364_inst_ack_1, ack => sendB_CP_2367_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: 	95 
    -- CP-element group 88: 	52 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/ptr_deref_1374_Split/$entry
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/ptr_deref_1374_Split/$exit
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/word_access_start/word_0/rr
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/word_access_start/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/word_access_start/$entry
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/ptr_deref_1374_Split/split_ack
      -- CP-element group 88: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/ptr_deref_1374_Split/split_req
      -- 
    rr_3297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(88), ack => ptr_deref_1374_store_0_req_0); -- 
    sendB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(87) & sendB_CP_2367_elements(95) & sendB_CP_2367_elements(52);
      gj_sendB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/word_access_start/word_0/ra
      -- CP-element group 89: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/word_access_start/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Sample/word_access_start/$exit
      -- 
    ra_3298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1374_store_0_ack_0, ack => sendB_CP_2367_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	52 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	96 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Update/word_access_complete/word_0/ca
      -- CP-element group 90: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Update/word_access_complete/word_0/$exit
      -- CP-element group 90: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Update/word_access_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1374_Update/$exit
      -- 
    ca_3309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1374_store_0_ack_1, ack => sendB_CP_2367_elements(90)); -- 
    -- CP-element group 91:  transition  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	64 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	68 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1269_ptr_deref_1290_delay
      -- 
    -- Element group sendB_CP_2367_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => sendB_CP_2367_elements(64), ack => sendB_CP_2367_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  transition  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	69 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	73 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1290_ptr_deref_1311_delay
      -- 
    -- Element group sendB_CP_2367_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => sendB_CP_2367_elements(69), ack => sendB_CP_2367_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  transition  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	74 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	78 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1311_ptr_deref_1332_delay
      -- 
    -- Element group sendB_CP_2367_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => sendB_CP_2367_elements(74), ack => sendB_CP_2367_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  transition  delay-element  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	79 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	83 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1332_ptr_deref_1353_delay
      -- 
    -- Element group sendB_CP_2367_elements(94) is a control-delay.
    cp_element_94_delay: control_delay_element  generic map(name => " 94_delay", delay_value => 1)  port map(req => sendB_CP_2367_elements(79), ack => sendB_CP_2367_elements(94), clk => clk, reset =>reset);
    -- CP-element group 95:  transition  delay-element  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	84 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	88 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/ptr_deref_1353_ptr_deref_1374_delay
      -- 
    -- Element group sendB_CP_2367_elements(95) is a control-delay.
    cp_element_95_delay: control_delay_element  generic map(name => " 95_delay", delay_value => 1)  port map(req => sendB_CP_2367_elements(84), ack => sendB_CP_2367_elements(95), clk => clk, reset =>reset);
    -- CP-element group 96:  branch  join  transition  place  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	85 
    -- CP-element group 96: 	90 
    -- CP-element group 96: 	54 
    -- CP-element group 96: 	55 
    -- CP-element group 96: 	75 
    -- CP-element group 96: 	80 
    -- CP-element group 96: 	70 
    -- CP-element group 96: 	65 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (10) 
      -- CP-element group 96: 	 branch_block_stmt_1002/R_cmp53x_xi_1384_place
      -- CP-element group 96: 	 branch_block_stmt_1002/if_stmt_1383_dead_link/$entry
      -- CP-element group 96: 	 branch_block_stmt_1002/if_stmt_1383_if_link/$entry
      -- CP-element group 96: 	 branch_block_stmt_1002/if_stmt_1383__entry__
      -- CP-element group 96: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382__exit__
      -- CP-element group 96: 	 branch_block_stmt_1002/if_stmt_1383_else_link/$entry
      -- CP-element group 96: 	 branch_block_stmt_1002/if_stmt_1383_eval_test/$exit
      -- CP-element group 96: 	 branch_block_stmt_1002/if_stmt_1383_eval_test/branch_req
      -- CP-element group 96: 	 branch_block_stmt_1002/assign_stmt_1239_to_assign_stmt_1382/$exit
      -- CP-element group 96: 	 branch_block_stmt_1002/if_stmt_1383_eval_test/$entry
      -- 
    branch_req_3322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(96), ack => if_stmt_1383_branch_req_0); -- 
    sendB_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(85) & sendB_CP_2367_elements(90) & sendB_CP_2367_elements(54) & sendB_CP_2367_elements(55) & sendB_CP_2367_elements(75) & sendB_CP_2367_elements(80) & sendB_CP_2367_elements(70) & sendB_CP_2367_elements(65);
      gj_sendB_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  place  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	137 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1002/ifx_xthen_sendRemainingElementsx_xexit
      -- CP-element group 97: 	 branch_block_stmt_1002/if_stmt_1383_if_link/if_choice_transition
      -- CP-element group 97: 	 branch_block_stmt_1002/if_stmt_1383_if_link/$exit
      -- CP-element group 97: 	 branch_block_stmt_1002/ifx_xthen_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 97: 	 branch_block_stmt_1002/ifx_xthen_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_3327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1383_branch_ack_1, ack => sendB_CP_2367_elements(97)); -- 
    -- CP-element group 98:  merge  transition  place  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	131 
    -- CP-element group 98:  members (18) 
      -- CP-element group 98: 	 branch_block_stmt_1002/if_stmt_1383_else_link/else_choice_transition
      -- CP-element group 98: 	 branch_block_stmt_1002/assign_stmt_1395_to_assign_stmt_1420__exit__
      -- CP-element group 98: 	 branch_block_stmt_1002/merge_stmt_1389__exit__
      -- CP-element group 98: 	 branch_block_stmt_1002/assign_stmt_1395_to_assign_stmt_1420__entry__
      -- CP-element group 98: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 98: 	 branch_block_stmt_1002/if_stmt_1383_else_link/$exit
      -- CP-element group 98: 	 branch_block_stmt_1002/ifx_xthen_bbx_xnphx_xi
      -- CP-element group 98: 	 branch_block_stmt_1002/assign_stmt_1395_to_assign_stmt_1420/$exit
      -- CP-element group 98: 	 branch_block_stmt_1002/assign_stmt_1395_to_assign_stmt_1420/$entry
      -- CP-element group 98: 	 branch_block_stmt_1002/ifx_xthen_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 98: 	 branch_block_stmt_1002/ifx_xthen_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 98: 	 branch_block_stmt_1002/merge_stmt_1389_PhiReqMerge
      -- CP-element group 98: 	 branch_block_stmt_1002/merge_stmt_1389_PhiAck/$entry
      -- CP-element group 98: 	 branch_block_stmt_1002/merge_stmt_1389_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_1002/merge_stmt_1389_PhiAck/dummy
      -- CP-element group 98: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 98: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/$entry
      -- CP-element group 98: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$entry
      -- 
    else_choice_transition_3331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1383_branch_ack_0, ack => sendB_CP_2367_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	136 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	116 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_sample_complete
      -- CP-element group 99: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_Sample/ack
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1441_index_offset_ack_0, ack => sendB_CP_2367_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	136 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (11) 
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_request/req
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_root_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_offset_calculated
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_request/$entry
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_base_plus_offset/sum_rename_ack
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_base_plus_offset/sum_rename_req
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_base_plus_offset/$exit
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_base_plus_offset/$entry
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_Update/ack
      -- CP-element group 100: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_Update/$exit
      -- 
    ack_3371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1441_index_offset_ack_1, ack => sendB_CP_2367_elements(100)); -- 
    req_3380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(100), ack => array_obj_ref_1441_final_reg_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_request/ack
      -- CP-element group 101: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_request/$exit
      -- 
    ack_3381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1441_final_reg_ack_0, ack => sendB_CP_2367_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	136 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	107 
    -- CP-element group 102:  members (24) 
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_complete/ack
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_word_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_root_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_address_resized
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_addr_resize/$entry
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_addr_resize/$exit
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_addr_resize/base_resize_req
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_addr_resize/base_resize_ack
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_plus_offset/$entry
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_plus_offset/$exit
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_plus_offset/sum_rename_req
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_base_plus_offset/sum_rename_ack
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_word_addrgen/$entry
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_word_addrgen/$exit
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_word_addrgen/root_register_req
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_word_addrgen/root_register_ack
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Sample/word_access_start/$entry
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Sample/word_access_start/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Sample/word_access_start/word_0/rr
      -- 
    ack_3386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1441_final_reg_ack_1, ack => sendB_CP_2367_elements(102)); -- 
    rr_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(102), ack => ptr_deref_1457_load_0_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	136 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	116 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_sample_complete
      -- CP-element group 103: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_Sample/ack
      -- 
    ack_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1453_index_offset_ack_0, ack => sendB_CP_2367_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	136 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (11) 
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_root_address_calculated
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_offset_calculated
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_base_plus_offset/$entry
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_base_plus_offset/$exit
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_base_plus_offset/sum_rename_req
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_base_plus_offset/sum_rename_ack
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_request/$entry
      -- CP-element group 104: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_request/req
      -- 
    ack_3418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1453_index_offset_ack_1, ack => sendB_CP_2367_elements(104)); -- 
    req_3427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(104), ack => array_obj_ref_1453_final_reg_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_request/$exit
      -- CP-element group 105: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_request/ack
      -- 
    ack_3428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1453_final_reg_ack_0, ack => sendB_CP_2367_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	136 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	111 
    -- CP-element group 106:  members (24) 
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_complete/$exit
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_complete/ack
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_word_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_root_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_address_resized
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_addr_resize/$entry
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_addr_resize/$exit
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_addr_resize/base_resize_req
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_addr_resize/base_resize_ack
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_plus_offset/$entry
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_plus_offset/$exit
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_plus_offset/sum_rename_req
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_base_plus_offset/sum_rename_ack
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_word_addrgen/$entry
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_word_addrgen/$exit
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_word_addrgen/root_register_req
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_word_addrgen/root_register_ack
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Sample/word_access_start/$entry
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Sample/word_access_start/word_0/$entry
      -- CP-element group 106: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Sample/word_access_start/word_0/rr
      -- 
    ack_3433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1453_final_reg_ack_1, ack => sendB_CP_2367_elements(106)); -- 
    rr_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(106), ack => ptr_deref_1464_load_0_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	102 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Sample/word_access_start/$exit
      -- CP-element group 107: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Sample/word_access_start/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Sample/word_access_start/word_0/ra
      -- 
    ra_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1457_load_0_ack_0, ack => sendB_CP_2367_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	136 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (12) 
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/word_access_complete/$exit
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/word_access_complete/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/word_access_complete/word_0/ca
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/ptr_deref_1457_Merge/$entry
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/ptr_deref_1457_Merge/$exit
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/ptr_deref_1457_Merge/merge_req
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/ptr_deref_1457_Merge/merge_ack
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_Sample/req
      -- 
    ca_3478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1457_load_0_ack_1, ack => sendB_CP_2367_elements(108)); -- 
    req_3491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(108), ack => WPIPE_maxpool_output_pipe_1459_inst_req_0); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_Sample/ack
      -- CP-element group 109: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_Update/req
      -- 
    ack_3492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1459_inst_ack_0, ack => sendB_CP_2367_elements(109)); -- 
    req_3496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(109), ack => WPIPE_maxpool_output_pipe_1459_inst_req_1); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1459_Update/ack
      -- 
    ack_3497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1459_inst_ack_1, ack => sendB_CP_2367_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	106 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Sample/word_access_start/$exit
      -- CP-element group 111: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Sample/word_access_start/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Sample/word_access_start/word_0/ra
      -- 
    ra_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1464_load_0_ack_0, ack => sendB_CP_2367_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	136 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/word_access_complete/$exit
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/word_access_complete/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/word_access_complete/word_0/ca
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/ptr_deref_1464_Merge/$entry
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/ptr_deref_1464_Merge/$exit
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/ptr_deref_1464_Merge/merge_req
      -- CP-element group 112: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/ptr_deref_1464_Merge/merge_ack
      -- 
    ca_3542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1464_load_0_ack_1, ack => sendB_CP_2367_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_Sample/req
      -- 
    req_3555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(113), ack => WPIPE_maxpool_output_pipe_1466_inst_req_0); -- 
    sendB_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(110) & sendB_CP_2367_elements(112);
      gj_sendB_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_update_start_
      -- CP-element group 114: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_Update/req
      -- 
    ack_3556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1466_inst_ack_0, ack => sendB_CP_2367_elements(114)); -- 
    req_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(114), ack => WPIPE_maxpool_output_pipe_1466_inst_req_1); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/WPIPE_maxpool_output_pipe_1466_Update/ack
      -- 
    ack_3561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1466_inst_ack_1, ack => sendB_CP_2367_elements(115)); -- 
    -- CP-element group 116:  branch  join  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: 	99 
    -- CP-element group 116: 	103 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_1002/if_stmt_1480__entry__
      -- CP-element group 116: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479__exit__
      -- CP-element group 116: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/$exit
      -- CP-element group 116: 	 branch_block_stmt_1002/if_stmt_1480_dead_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_1002/if_stmt_1480_eval_test/$entry
      -- CP-element group 116: 	 branch_block_stmt_1002/if_stmt_1480_eval_test/$exit
      -- CP-element group 116: 	 branch_block_stmt_1002/if_stmt_1480_eval_test/branch_req
      -- CP-element group 116: 	 branch_block_stmt_1002/R_exitcond1_1481_place
      -- CP-element group 116: 	 branch_block_stmt_1002/if_stmt_1480_if_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_1002/if_stmt_1480_else_link/$entry
      -- 
    branch_req_3569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(116), ack => if_stmt_1480_branch_req_0); -- 
    sendB_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(115) & sendB_CP_2367_elements(99) & sendB_CP_2367_elements(103);
      gj_sendB_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  merge  transition  place  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	137 
    -- CP-element group 117:  members (13) 
      -- CP-element group 117: 	 branch_block_stmt_1002/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit
      -- CP-element group 117: 	 branch_block_stmt_1002/merge_stmt_1486__exit__
      -- CP-element group 117: 	 branch_block_stmt_1002/if_stmt_1480_if_link/$exit
      -- CP-element group 117: 	 branch_block_stmt_1002/if_stmt_1480_if_link/if_choice_transition
      -- CP-element group 117: 	 branch_block_stmt_1002/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit
      -- CP-element group 117: 	 branch_block_stmt_1002/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 117: 	 branch_block_stmt_1002/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit_PhiReq/$exit
      -- CP-element group 117: 	 branch_block_stmt_1002/merge_stmt_1486_PhiReqMerge
      -- CP-element group 117: 	 branch_block_stmt_1002/merge_stmt_1486_PhiAck/$entry
      -- CP-element group 117: 	 branch_block_stmt_1002/merge_stmt_1486_PhiAck/$exit
      -- CP-element group 117: 	 branch_block_stmt_1002/merge_stmt_1486_PhiAck/dummy
      -- CP-element group 117: 	 branch_block_stmt_1002/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 117: 	 branch_block_stmt_1002/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_3574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1480_branch_ack_1, ack => sendB_CP_2367_elements(117)); -- 
    -- CP-element group 118:  fork  transition  place  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	132 
    -- CP-element group 118: 	133 
    -- CP-element group 118:  members (12) 
      -- CP-element group 118: 	 branch_block_stmt_1002/if_stmt_1480_else_link/$exit
      -- CP-element group 118: 	 branch_block_stmt_1002/if_stmt_1480_else_link/else_choice_transition
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/$entry
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$entry
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/$entry
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/$entry
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1480_branch_ack_0, ack => sendB_CP_2367_elements(118)); -- 
    rr_3742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(118), ack => type_cast_1429_inst_req_0); -- 
    cr_3747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(118), ack => type_cast_1429_inst_req_1); -- 
    -- CP-element group 119:  transition  output  delay-element  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	1 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1049/$exit
      -- CP-element group 119: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1053_konst_delay_trans
      -- CP-element group 119: 	 branch_block_stmt_1002/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_req
      -- 
    phi_stmt_1049_req_3603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1049_req_3603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(119), ack => phi_stmt_1049_req_0); -- 
    -- Element group sendB_CP_2367_elements(119) is a control-delay.
    cp_element_119_delay: control_delay_element  generic map(name => " 119_delay", delay_value => 1)  port map(req => sendB_CP_2367_elements(1), ack => sendB_CP_2367_elements(119), clk => clk, reset =>reset);
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	50 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/Sample/ra
      -- 
    ra_3623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_0, ack => sendB_CP_2367_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	50 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/Update/ca
      -- 
    ca_3628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_1, ack => sendB_CP_2367_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (6) 
      -- CP-element group 122: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/$exit
      -- CP-element group 122: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/$exit
      -- CP-element group 122: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_sources/type_cast_1055/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_1002/forx_xbody_forx_xbody_PhiReq/phi_stmt_1049/phi_stmt_1049_req
      -- 
    phi_stmt_1049_req_3629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1049_req_3629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(122), ack => phi_stmt_1049_req_1); -- 
    sendB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(120) & sendB_CP_2367_elements(121);
      gj_sendB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1002/merge_stmt_1048_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_1002/merge_stmt_1048_PhiAck/$entry
      -- 
    sendB_CP_2367_elements(123) <= OrReduce(sendB_CP_2367_elements(119) & sendB_CP_2367_elements(122));
    -- CP-element group 124:  fork  transition  place  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: 	16 
    -- CP-element group 124: 	18 
    -- CP-element group 124: 	20 
    -- CP-element group 124: 	22 
    -- CP-element group 124: 	24 
    -- CP-element group 124: 	3 
    -- CP-element group 124: 	4 
    -- CP-element group 124: 	6 
    -- CP-element group 124: 	10 
    -- CP-element group 124: 	12 
    -- CP-element group 124: 	14 
    -- CP-element group 124:  members (53) 
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_scaled_1
      -- CP-element group 124: 	 branch_block_stmt_1002/merge_stmt_1048__exit__
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/word_access_complete/word_0/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_computed_1
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_resize_1/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_resize_1/$exit
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176__entry__
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_resize_1/index_resize_req
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1080_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_resize_1/index_resize_ack
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1070_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_resized_1
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_complete/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_scale_1/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_scale_1/$exit
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/addr_of_1062_complete/req
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_update_start
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/word_access_complete/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_Update/req
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_final_index_sum_regn_Sample/req
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/ptr_deref_1066_Update/word_access_complete/word_0/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_scale_1/scale_rename_ack
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/array_obj_ref_1061_index_scale_1/scale_rename_req
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1090_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1100_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1110_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1120_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1130_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_update_start_
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1002/assign_stmt_1063_to_assign_stmt_1176/type_cast_1140_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_1002/merge_stmt_1048_PhiAck/$exit
      -- CP-element group 124: 	 branch_block_stmt_1002/merge_stmt_1048_PhiAck/phi_stmt_1049_ack
      -- 
    phi_stmt_1049_ack_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1049_ack_0, ack => sendB_CP_2367_elements(124)); -- 
    cr_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => ptr_deref_1066_load_0_req_1); -- 
    cr_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => type_cast_1080_inst_req_1); -- 
    cr_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => type_cast_1070_inst_req_1); -- 
    req_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => addr_of_1062_final_reg_req_1); -- 
    req_2478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => array_obj_ref_1061_index_offset_req_1); -- 
    req_2473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => array_obj_ref_1061_index_offset_req_0); -- 
    cr_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => type_cast_1090_inst_req_1); -- 
    cr_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => type_cast_1100_inst_req_1); -- 
    cr_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => type_cast_1110_inst_req_1); -- 
    cr_2627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => type_cast_1120_inst_req_1); -- 
    cr_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => type_cast_1130_inst_req_1); -- 
    cr_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(124), ack => type_cast_1140_inst_req_1); -- 
    -- CP-element group 125:  transition  output  delay-element  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	2 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1002/entry_forx_xend_PhiReq/$exit
      -- CP-element group 125: 	 branch_block_stmt_1002/entry_forx_xend_PhiReq/phi_stmt_1209/$exit
      -- CP-element group 125: 	 branch_block_stmt_1002/entry_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_1002/entry_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1215_konst_delay_trans
      -- CP-element group 125: 	 branch_block_stmt_1002/entry_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_req
      -- 
    phi_stmt_1209_req_3657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1209_req_3657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(125), ack => phi_stmt_1209_req_1); -- 
    -- Element group sendB_CP_2367_elements(125) is a control-delay.
    cp_element_125_delay: control_delay_element  generic map(name => " 125_delay", delay_value => 1)  port map(req => sendB_CP_2367_elements(2), ack => sendB_CP_2367_elements(125), clk => clk, reset =>reset);
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	49 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/Sample/ra
      -- 
    ra_3677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1212_inst_ack_0, ack => sendB_CP_2367_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	49 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/Update/ca
      -- 
    ca_3682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1212_inst_ack_1, ack => sendB_CP_2367_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 128: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/$exit
      -- CP-element group 128: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/$exit
      -- CP-element group 128: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_sources/type_cast_1212/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_1002/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1209/phi_stmt_1209_req
      -- 
    phi_stmt_1209_req_3683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1209_req_3683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(128), ack => phi_stmt_1209_req_0); -- 
    sendB_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(126) & sendB_CP_2367_elements(127);
      gj_sendB_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  merge  transition  place  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	125 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_1002/merge_stmt_1208_PhiReqMerge
      -- CP-element group 129: 	 branch_block_stmt_1002/merge_stmt_1208_PhiAck/$entry
      -- 
    sendB_CP_2367_elements(129) <= OrReduce(sendB_CP_2367_elements(125) & sendB_CP_2367_elements(128));
    -- CP-element group 130:  branch  transition  place  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	51 
    -- CP-element group 130: 	52 
    -- CP-element group 130:  members (15) 
      -- CP-element group 130: 	 branch_block_stmt_1002/merge_stmt_1208__exit__
      -- CP-element group 130: 	 branch_block_stmt_1002/assign_stmt_1222_to_assign_stmt_1228__entry__
      -- CP-element group 130: 	 branch_block_stmt_1002/assign_stmt_1222_to_assign_stmt_1228__exit__
      -- CP-element group 130: 	 branch_block_stmt_1002/if_stmt_1229__entry__
      -- CP-element group 130: 	 branch_block_stmt_1002/assign_stmt_1222_to_assign_stmt_1228/$entry
      -- CP-element group 130: 	 branch_block_stmt_1002/assign_stmt_1222_to_assign_stmt_1228/$exit
      -- CP-element group 130: 	 branch_block_stmt_1002/if_stmt_1229_dead_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_1002/if_stmt_1229_eval_test/$entry
      -- CP-element group 130: 	 branch_block_stmt_1002/if_stmt_1229_eval_test/$exit
      -- CP-element group 130: 	 branch_block_stmt_1002/if_stmt_1229_eval_test/branch_req
      -- CP-element group 130: 	 branch_block_stmt_1002/R_tobool_1230_place
      -- CP-element group 130: 	 branch_block_stmt_1002/if_stmt_1229_if_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_1002/if_stmt_1229_else_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_1002/merge_stmt_1208_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_1002/merge_stmt_1208_PhiAck/phi_stmt_1209_ack
      -- 
    phi_stmt_1209_ack_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1209_ack_0, ack => sendB_CP_2367_elements(130)); -- 
    branch_req_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(130), ack => if_stmt_1229_branch_req_0); -- 
    -- CP-element group 131:  transition  output  delay-element  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	98 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	135 
    -- CP-element group 131:  members (5) 
      -- CP-element group 131: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- CP-element group 131: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/$exit
      -- CP-element group 131: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$exit
      -- CP-element group 131: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1427_konst_delay_trans
      -- CP-element group 131: 	 branch_block_stmt_1002/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_req
      -- 
    phi_stmt_1423_req_3723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1423_req_3723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(131), ack => phi_stmt_1423_req_0); -- 
    -- Element group sendB_CP_2367_elements(131) is a control-delay.
    cp_element_131_delay: control_delay_element  generic map(name => " 131_delay", delay_value => 1)  port map(req => sendB_CP_2367_elements(98), ack => sendB_CP_2367_elements(131), clk => clk, reset =>reset);
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	118 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/ra
      -- 
    ra_3743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_0, ack => sendB_CP_2367_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	118 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (2) 
      -- CP-element group 133: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/ca
      -- 
    ca_3748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_1, ack => sendB_CP_2367_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- CP-element group 134: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/$exit
      -- CP-element group 134: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$exit
      -- CP-element group 134: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/$exit
      -- CP-element group 134: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/$exit
      -- CP-element group 134: 	 branch_block_stmt_1002/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1423/phi_stmt_1423_req
      -- 
    phi_stmt_1423_req_3749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1423_req_3749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(134), ack => phi_stmt_1423_req_1); -- 
    sendB_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2367_elements(132) & sendB_CP_2367_elements(133);
      gj_sendB_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2367_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  merge  transition  place  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	131 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_1002/merge_stmt_1422_PhiReqMerge
      -- CP-element group 135: 	 branch_block_stmt_1002/merge_stmt_1422_PhiAck/$entry
      -- 
    sendB_CP_2367_elements(135) <= OrReduce(sendB_CP_2367_elements(131) & sendB_CP_2367_elements(134));
    -- CP-element group 136:  fork  transition  place  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	108 
    -- CP-element group 136: 	112 
    -- CP-element group 136: 	99 
    -- CP-element group 136: 	100 
    -- CP-element group 136: 	102 
    -- CP-element group 136: 	103 
    -- CP-element group 136: 	104 
    -- CP-element group 136: 	106 
    -- CP-element group 136:  members (53) 
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_resize_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_resize_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_computed_1
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_scaled_1
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_resize_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_resize_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_resized_1
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_computed_1
      -- CP-element group 136: 	 branch_block_stmt_1002/merge_stmt_1422__exit__
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479__entry__
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_scaled_1
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_resize_1/index_resize_req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_resize_1/index_resize_ack
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_resize_1/index_resize_req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_scale_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_scale_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_scale_1/scale_rename_req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_scale_1/scale_rename_ack
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_update_start_
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_index_resized_1
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_complete/req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_update_start_
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_update_start
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_Update/req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_Sample/req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1441_final_index_sum_regn_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_resize_1/index_resize_ack
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_scale_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_scale_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_scale_1/scale_rename_req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_index_scale_1/scale_rename_ack
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_update_start
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_Sample/req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_final_index_sum_regn_Update/req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/array_obj_ref_1453_complete/req
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_update_start_
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/word_access_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/word_access_complete/word_0/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1457_Update/word_access_complete/word_0/cr
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_update_start_
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/word_access_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/word_access_complete/word_0/$entry
      -- CP-element group 136: 	 branch_block_stmt_1002/assign_stmt_1436_to_assign_stmt_1479/ptr_deref_1464_Update/word_access_complete/word_0/cr
      -- CP-element group 136: 	 branch_block_stmt_1002/merge_stmt_1422_PhiAck/$exit
      -- CP-element group 136: 	 branch_block_stmt_1002/merge_stmt_1422_PhiAck/phi_stmt_1423_ack
      -- 
    phi_stmt_1423_ack_3754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1423_ack_0, ack => sendB_CP_2367_elements(136)); -- 
    req_3385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(136), ack => array_obj_ref_1441_final_reg_req_1); -- 
    req_3370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(136), ack => array_obj_ref_1441_index_offset_req_1); -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(136), ack => array_obj_ref_1441_index_offset_req_0); -- 
    req_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(136), ack => array_obj_ref_1453_index_offset_req_0); -- 
    req_3417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(136), ack => array_obj_ref_1453_index_offset_req_1); -- 
    req_3432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(136), ack => array_obj_ref_1453_final_reg_req_1); -- 
    cr_3477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(136), ack => ptr_deref_1457_load_0_req_1); -- 
    cr_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2367_elements(136), ack => ptr_deref_1464_load_0_req_1); -- 
    -- CP-element group 137:  merge  transition  place  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	117 
    -- CP-element group 137: 	97 
    -- CP-element group 137: 	51 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (16) 
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1490__exit__
      -- CP-element group 137: 	 branch_block_stmt_1002/return__
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1488__exit__
      -- CP-element group 137: 	 branch_block_stmt_1002/branch_block_stmt_1002__exit__
      -- CP-element group 137: 	 branch_block_stmt_1002/$exit
      -- CP-element group 137: 	 $exit
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1490_PhiReqMerge
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1488_PhiReqMerge
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1488_PhiAck/$entry
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1488_PhiAck/$exit
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1488_PhiAck/dummy
      -- CP-element group 137: 	 branch_block_stmt_1002/return___PhiReq/$entry
      -- CP-element group 137: 	 branch_block_stmt_1002/return___PhiReq/$exit
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1490_PhiAck/$entry
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1490_PhiAck/$exit
      -- CP-element group 137: 	 branch_block_stmt_1002/merge_stmt_1490_PhiAck/dummy
      -- 
    sendB_CP_2367_elements(137) <= OrReduce(sendB_CP_2367_elements(117) & sendB_CP_2367_elements(97) & sendB_CP_2367_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1204_wire : std_logic_vector(63 downto 0);
    signal R_indvar_1060_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1060_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1243_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1243_scaled : std_logic_vector(13 downto 0);
    signal R_tmp2_1440_resized : std_logic_vector(2 downto 0);
    signal R_tmp2_1440_scaled : std_logic_vector(2 downto 0);
    signal R_tmp3_1452_resized : std_logic_vector(2 downto 0);
    signal R_tmp3_1452_scaled : std_logic_vector(2 downto 0);
    signal and70_1222 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1061_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1061_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1061_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1061_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1061_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1061_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1441_constant_part_of_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1441_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1441_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1441_offset_scale_factor_1 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1441_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1441_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1453_constant_part_of_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1453_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1453_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1453_offset_scale_factor_1 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1453_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1453_root_address : std_logic_vector(2 downto 0);
    signal arrayidx11x_xi_1288 : std_logic_vector(31 downto 0);
    signal arrayidx17x_xi_1309 : std_logic_vector(31 downto 0);
    signal arrayidx23x_xi_1330 : std_logic_vector(31 downto 0);
    signal arrayidx29x_xi_1351 : std_logic_vector(31 downto 0);
    signal arrayidx35x_xi_1372 : std_logic_vector(31 downto 0);
    signal arrayidx43x_xi_1442 : std_logic_vector(31 downto 0);
    signal arrayidx48x_xi_1454 : std_logic_vector(31 downto 0);
    signal arrayidx5x_xi_1267 : std_logic_vector(31 downto 0);
    signal arrayidx_1063 : std_logic_vector(31 downto 0);
    signal arrayidxx_xi_1246 : std_logic_vector(31 downto 0);
    signal cmp53x_xi_1382 : std_logic_vector(0 downto 0);
    signal cmp77_1014 : std_logic_vector(0 downto 0);
    signal conv10x_xi_1281 : std_logic_vector(7 downto 0);
    signal conv14_1081 : std_logic_vector(7 downto 0);
    signal conv16x_xi_1302 : std_logic_vector(7 downto 0);
    signal conv20_1091 : std_logic_vector(7 downto 0);
    signal conv22x_xi_1323 : std_logic_vector(7 downto 0);
    signal conv26_1101 : std_logic_vector(7 downto 0);
    signal conv28x_xi_1344 : std_logic_vector(7 downto 0);
    signal conv32_1111 : std_logic_vector(7 downto 0);
    signal conv34x_xi_1365 : std_logic_vector(7 downto 0);
    signal conv38_1121 : std_logic_vector(7 downto 0);
    signal conv44_1131 : std_logic_vector(7 downto 0);
    signal conv50_1141 : std_logic_vector(7 downto 0);
    signal conv74_1239 : std_logic_vector(15 downto 0);
    signal conv8_1071 : std_logic_vector(7 downto 0);
    signal convx_xi_1260 : std_logic_vector(7 downto 0);
    signal exitcond1_1479 : std_logic_vector(0 downto 0);
    signal exitcond_1176 : std_logic_vector(0 downto 0);
    signal iNsTr_29_1407 : std_logic_vector(63 downto 0);
    signal indvar_1049 : std_logic_vector(63 downto 0);
    signal indvarx_xi_1423 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1171 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi_1474 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_1209 : std_logic_vector(63 downto 0);
    signal out_datax_xi_1008 : std_logic_vector(31 downto 0);
    signal phitmp_1206 : std_logic_vector(63 downto 0);
    signal ptr_deref_1066_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1066_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1066_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1066_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1066_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1249_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1249_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1249_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1249_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1249_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1269_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1269_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1269_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1269_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1269_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1269_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1290_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1290_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1290_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1290_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1290_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1290_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1311_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1311_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1311_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1311_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1311_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1311_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1332_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1332_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1332_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1332_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1332_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1332_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1353_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1353_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1353_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1353_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1353_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1353_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1374_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1374_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1374_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1374_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1374_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1374_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1457_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1457_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1457_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1457_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1457_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1464_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1464_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1464_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1464_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1464_word_offset_0 : std_logic_vector(2 downto 0);
    signal shr11_1077 : std_logic_vector(63 downto 0);
    signal shr13x_xi_1298 : std_logic_vector(63 downto 0);
    signal shr17_1087 : std_logic_vector(63 downto 0);
    signal shr19x_xi_1319 : std_logic_vector(63 downto 0);
    signal shr23_1097 : std_logic_vector(63 downto 0);
    signal shr25x_xi_1340 : std_logic_vector(63 downto 0);
    signal shr29_1107 : std_logic_vector(63 downto 0);
    signal shr31x_xi_1361 : std_logic_vector(63 downto 0);
    signal shr35_1117 : std_logic_vector(63 downto 0);
    signal shr41_1127 : std_logic_vector(63 downto 0);
    signal shr47_1137 : std_logic_vector(63 downto 0);
    signal shr7x_xi_1277 : std_logic_vector(63 downto 0);
    signal shr_1027 : std_logic_vector(63 downto 0);
    signal shrx_xi_1256 : std_logic_vector(63 downto 0);
    signal tmp1x_xi_1250 : std_logic_vector(63 downto 0);
    signal tmp2_1436 : std_logic_vector(63 downto 0);
    signal tmp3_1448 : std_logic_vector(63 downto 0);
    signal tmp44x_xi_1458 : std_logic_vector(7 downto 0);
    signal tmp49x_xi_1465 : std_logic_vector(7 downto 0);
    signal tmp55x_xi_1395 : std_logic_vector(0 downto 0);
    signal tmp58x_xi_1420 : std_logic_vector(63 downto 0);
    signal tmp5_1067 : std_logic_vector(63 downto 0);
    signal tmp80_1033 : std_logic_vector(0 downto 0);
    signal tmp81_1196 : std_logic_vector(63 downto 0);
    signal tmp_1039 : std_logic_vector(0 downto 0);
    signal tmpx_xopx_xi_1401 : std_logic_vector(63 downto 0);
    signal tobool_1228 : std_logic_vector(0 downto 0);
    signal type_cast_1012_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1025_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1031_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1037_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1044_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1053_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1055_wire : std_logic_vector(63 downto 0);
    signal type_cast_1075_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1085_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1095_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1105_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1115_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1125_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1135_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1169_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1188_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1194_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1200_wire : std_logic_vector(63 downto 0);
    signal type_cast_1203_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1212_wire : std_logic_vector(63 downto 0);
    signal type_cast_1215_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1220_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1226_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1275_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1296_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1317_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1359_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1380_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1393_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1399_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1405_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1411_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1418_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1427_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1429_wire : std_logic_vector(63 downto 0);
    signal type_cast_1434_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1446_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1472_wire_constant : std_logic_vector(63 downto 0);
    signal umax4_1046 : std_logic_vector(63 downto 0);
    signal umax_1190 : std_logic_vector(63 downto 0);
    signal xx_xopx_xi_1413 : std_logic_vector(63 downto 0);
    signal xxsendBxxbodyxxout_datax_xi_alloc_base_address : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    array_obj_ref_1061_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1061_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1061_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1061_resized_base_address <= "00000000000000";
    array_obj_ref_1244_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1244_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1244_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1244_resized_base_address <= "00000000000000";
    array_obj_ref_1441_constant_part_of_offset <= "000";
    array_obj_ref_1441_offset_scale_factor_0 <= "110";
    array_obj_ref_1441_offset_scale_factor_1 <= "001";
    array_obj_ref_1441_resized_base_address <= "000";
    array_obj_ref_1453_constant_part_of_offset <= "000";
    array_obj_ref_1453_offset_scale_factor_0 <= "110";
    array_obj_ref_1453_offset_scale_factor_1 <= "001";
    array_obj_ref_1453_resized_base_address <= "000";
    arrayidx11x_xi_1288 <= "00000000000000000000000000000100";
    arrayidx17x_xi_1309 <= "00000000000000000000000000000011";
    arrayidx23x_xi_1330 <= "00000000000000000000000000000010";
    arrayidx29x_xi_1351 <= "00000000000000000000000000000001";
    arrayidx35x_xi_1372 <= "00000000000000000000000000000000";
    arrayidx5x_xi_1267 <= "00000000000000000000000000000101";
    out_datax_xi_1008 <= "00000000000000000000000000000000";
    ptr_deref_1066_word_offset_0 <= "00000000000000";
    ptr_deref_1249_word_offset_0 <= "00000000000000";
    ptr_deref_1269_word_offset_0 <= "000";
    ptr_deref_1290_word_offset_0 <= "000";
    ptr_deref_1311_word_offset_0 <= "000";
    ptr_deref_1332_word_offset_0 <= "000";
    ptr_deref_1353_word_offset_0 <= "000";
    ptr_deref_1374_word_offset_0 <= "000";
    ptr_deref_1457_word_offset_0 <= "000";
    ptr_deref_1464_word_offset_0 <= "000";
    type_cast_1012_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1025_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1031_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1037_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1044_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1053_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1075_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1085_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1095_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1105_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1115_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1125_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1135_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1169_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1188_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1194_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1203_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1215_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1220_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1226_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1254_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1275_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1296_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1317_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1338_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1359_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1380_wire_constant <= "0000000000000000";
    type_cast_1393_wire_constant <= "0000000000000001";
    type_cast_1399_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_1405_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_1411_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1418_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1427_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1434_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1446_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1472_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    xxsendBxxbodyxxout_datax_xi_alloc_base_address <= "000";
    phi_stmt_1049: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1053_wire_constant & type_cast_1055_wire;
      req <= phi_stmt_1049_req_0 & phi_stmt_1049_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1049",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1049_ack_0,
          idata => idata,
          odata => indvar_1049,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1049
    phi_stmt_1209: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1212_wire & type_cast_1215_wire_constant;
      req <= phi_stmt_1209_req_0 & phi_stmt_1209_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1209",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1209_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_1209,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1209
    phi_stmt_1423: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1427_wire_constant & type_cast_1429_wire;
      req <= phi_stmt_1423_req_0 & phi_stmt_1423_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1423",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1423_ack_0,
          idata => idata,
          odata => indvarx_xi_1423,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1423
    -- flow-through select operator MUX_1045_inst
    umax4_1046 <= shr_1027 when (tmp_1039(0) /=  '0') else type_cast_1044_wire_constant;
    -- flow-through select operator MUX_1189_inst
    umax_1190 <= shr_1027 when (tmp80_1033(0) /=  '0') else type_cast_1188_wire_constant;
    -- flow-through select operator MUX_1419_inst
    tmp58x_xi_1420 <= xx_xopx_xi_1413 when (tmp55x_xi_1395(0) /=  '0') else type_cast_1418_wire_constant;
    addr_of_1062_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1062_final_reg_req_0;
      addr_of_1062_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1062_final_reg_req_1;
      addr_of_1062_final_reg_ack_1<= rack(0);
      addr_of_1062_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1062_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1061_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1063,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1245_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1245_final_reg_req_0;
      addr_of_1245_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1245_final_reg_req_1;
      addr_of_1245_final_reg_ack_1<= rack(0);
      addr_of_1245_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1245_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1244_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidxx_xi_1246,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    array_obj_ref_1441_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= array_obj_ref_1441_final_reg_req_0;
      array_obj_ref_1441_final_reg_ack_0<= wack(0);
      rreq(0) <= array_obj_ref_1441_final_reg_req_1;
      array_obj_ref_1441_final_reg_ack_1<= rack(0);
      array_obj_ref_1441_final_reg : InterlockBuffer generic map ( -- 
        name => "array_obj_ref_1441_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1441_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx43x_xi_1442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    array_obj_ref_1453_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= array_obj_ref_1453_final_reg_req_0;
      array_obj_ref_1453_final_reg_ack_0<= wack(0);
      rreq(0) <= array_obj_ref_1453_final_reg_req_1;
      array_obj_ref_1453_final_reg_ack_1<= rack(0);
      array_obj_ref_1453_final_reg : InterlockBuffer generic map ( -- 
        name => "array_obj_ref_1453_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1453_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx48x_xi_1454,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1055_inst_req_0;
      type_cast_1055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1055_inst_req_1;
      type_cast_1055_inst_ack_1<= rack(0);
      type_cast_1055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1055_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1070_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1070_inst_req_0;
      type_cast_1070_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1070_inst_req_1;
      type_cast_1070_inst_ack_1<= rack(0);
      type_cast_1070_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1070_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_1067,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_1071,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1080_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1080_inst_req_0;
      type_cast_1080_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1080_inst_req_1;
      type_cast_1080_inst_ack_1<= rack(0);
      type_cast_1080_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1080_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr11_1077,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_1081,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1090_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1090_inst_req_0;
      type_cast_1090_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1090_inst_req_1;
      type_cast_1090_inst_ack_1<= rack(0);
      type_cast_1090_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1090_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_1087,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_1091,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1100_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1100_inst_req_0;
      type_cast_1100_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1100_inst_req_1;
      type_cast_1100_inst_ack_1<= rack(0);
      type_cast_1100_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1100_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_1097,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_1101,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1110_inst_req_0;
      type_cast_1110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1110_inst_req_1;
      type_cast_1110_inst_ack_1<= rack(0);
      type_cast_1110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_1107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1120_inst_req_0;
      type_cast_1120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1120_inst_req_1;
      type_cast_1120_inst_ack_1<= rack(0);
      type_cast_1120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_1117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_1121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1130_inst_req_0;
      type_cast_1130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1130_inst_req_1;
      type_cast_1130_inst_ack_1<= rack(0);
      type_cast_1130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_1127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_1131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1140_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1140_inst_req_0;
      type_cast_1140_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1140_inst_req_1;
      type_cast_1140_inst_ack_1<= rack(0);
      type_cast_1140_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1140_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr47_1137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_1141,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1200_inst
    process(tmp81_1196) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp81_1196(63 downto 0);
      type_cast_1200_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1205_inst
    process(ASHR_i64_i64_1204_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1204_wire(63 downto 0);
      phitmp_1206 <= tmp_var; -- 
    end process;
    type_cast_1212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1212_inst_req_0;
      type_cast_1212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1212_inst_req_1;
      type_cast_1212_inst_ack_1<= rack(0);
      type_cast_1212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_1206,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1212_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => and70_1222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1259_inst_req_0;
      type_cast_1259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1259_inst_req_1;
      type_cast_1259_inst_ack_1<= rack(0);
      type_cast_1259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xi_1256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1280_inst_req_0;
      type_cast_1280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1280_inst_req_1;
      type_cast_1280_inst_ack_1<= rack(0);
      type_cast_1280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr7x_xi_1277,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10x_xi_1281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1301_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1301_inst_req_0;
      type_cast_1301_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1301_inst_req_1;
      type_cast_1301_inst_ack_1<= rack(0);
      type_cast_1301_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1301_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr13x_xi_1298,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16x_xi_1302,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1322_inst_req_0;
      type_cast_1322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1322_inst_req_1;
      type_cast_1322_inst_ack_1<= rack(0);
      type_cast_1322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr19x_xi_1319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22x_xi_1323,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1343_inst_req_0;
      type_cast_1343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1343_inst_req_1;
      type_cast_1343_inst_ack_1<= rack(0);
      type_cast_1343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr25x_xi_1340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28x_xi_1344,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1364_inst_req_0;
      type_cast_1364_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1364_inst_req_1;
      type_cast_1364_inst_ack_1<= rack(0);
      type_cast_1364_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1364_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr31x_xi_1361,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34x_xi_1365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1429_inst_req_0;
      type_cast_1429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1429_inst_req_1;
      type_cast_1429_inst_ack_1<= rack(0);
      type_cast_1429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi_1474,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1429_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1061_index_1_rename
    process(R_indvar_1060_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1060_resized;
      ov(13 downto 0) := iv;
      R_indvar_1060_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1061_index_1_resize
    process(indvar_1049) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1049;
      ov := iv(13 downto 0);
      R_indvar_1060_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1061_root_address_inst
    process(array_obj_ref_1061_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1061_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1061_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1244_index_1_rename
    process(R_ix_x0x_xlcssa_1243_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1243_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1243_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1244_index_1_resize
    process(ix_x0x_xlcssa_1209) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_1209;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1243_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1244_root_address_inst
    process(array_obj_ref_1244_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1244_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1244_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_index_1_rename
    process(R_tmp2_1440_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp2_1440_resized;
      ov(2 downto 0) := iv;
      R_tmp2_1440_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_index_1_resize
    process(tmp2_1436) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp2_1436;
      ov := iv(2 downto 0);
      R_tmp2_1440_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_root_address_inst
    process(array_obj_ref_1441_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1441_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_1441_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1453_index_1_rename
    process(R_tmp3_1452_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp3_1452_resized;
      ov(2 downto 0) := iv;
      R_tmp3_1452_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1453_index_1_resize
    process(tmp3_1448) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp3_1448;
      ov := iv(2 downto 0);
      R_tmp3_1452_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1453_root_address_inst
    process(array_obj_ref_1453_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1453_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_1453_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1066_addr_0
    process(ptr_deref_1066_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1066_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1066_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1066_base_resize
    process(arrayidx_1063) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1063;
      ov := iv(13 downto 0);
      ptr_deref_1066_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1066_gather_scatter
    process(ptr_deref_1066_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1066_data_0;
      ov(63 downto 0) := iv;
      tmp5_1067 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1066_root_address_inst
    process(ptr_deref_1066_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1066_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1066_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1249_addr_0
    process(ptr_deref_1249_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1249_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1249_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1249_base_resize
    process(arrayidxx_xi_1246) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidxx_xi_1246;
      ov := iv(13 downto 0);
      ptr_deref_1249_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1249_gather_scatter
    process(ptr_deref_1249_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1249_data_0;
      ov(63 downto 0) := iv;
      tmp1x_xi_1250 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1249_root_address_inst
    process(ptr_deref_1249_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1249_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1249_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1269_addr_0
    process(ptr_deref_1269_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1269_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1269_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1269_base_resize
    process(arrayidx5x_xi_1267) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx5x_xi_1267;
      ov := iv(2 downto 0);
      ptr_deref_1269_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1269_gather_scatter
    process(convx_xi_1260) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := convx_xi_1260;
      ov(7 downto 0) := iv;
      ptr_deref_1269_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1269_root_address_inst
    process(ptr_deref_1269_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1269_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1269_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1290_addr_0
    process(ptr_deref_1290_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1290_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1290_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1290_base_resize
    process(arrayidx11x_xi_1288) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx11x_xi_1288;
      ov := iv(2 downto 0);
      ptr_deref_1290_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1290_gather_scatter
    process(conv10x_xi_1281) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv10x_xi_1281;
      ov(7 downto 0) := iv;
      ptr_deref_1290_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1290_root_address_inst
    process(ptr_deref_1290_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1290_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1290_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1311_addr_0
    process(ptr_deref_1311_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1311_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1311_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1311_base_resize
    process(arrayidx17x_xi_1309) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx17x_xi_1309;
      ov := iv(2 downto 0);
      ptr_deref_1311_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1311_gather_scatter
    process(conv16x_xi_1302) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv16x_xi_1302;
      ov(7 downto 0) := iv;
      ptr_deref_1311_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1311_root_address_inst
    process(ptr_deref_1311_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1311_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1311_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1332_addr_0
    process(ptr_deref_1332_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1332_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1332_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1332_base_resize
    process(arrayidx23x_xi_1330) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx23x_xi_1330;
      ov := iv(2 downto 0);
      ptr_deref_1332_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1332_gather_scatter
    process(conv22x_xi_1323) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv22x_xi_1323;
      ov(7 downto 0) := iv;
      ptr_deref_1332_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1332_root_address_inst
    process(ptr_deref_1332_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1332_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1332_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1353_addr_0
    process(ptr_deref_1353_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1353_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1353_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1353_base_resize
    process(arrayidx29x_xi_1351) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx29x_xi_1351;
      ov := iv(2 downto 0);
      ptr_deref_1353_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1353_gather_scatter
    process(conv28x_xi_1344) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv28x_xi_1344;
      ov(7 downto 0) := iv;
      ptr_deref_1353_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1353_root_address_inst
    process(ptr_deref_1353_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1353_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1353_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1374_addr_0
    process(ptr_deref_1374_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1374_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1374_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1374_base_resize
    process(arrayidx35x_xi_1372) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx35x_xi_1372;
      ov := iv(2 downto 0);
      ptr_deref_1374_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1374_gather_scatter
    process(conv34x_xi_1365) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv34x_xi_1365;
      ov(7 downto 0) := iv;
      ptr_deref_1374_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1374_root_address_inst
    process(ptr_deref_1374_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1374_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1374_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1457_addr_0
    process(ptr_deref_1457_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1457_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1457_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1457_base_resize
    process(arrayidx43x_xi_1442) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx43x_xi_1442;
      ov := iv(2 downto 0);
      ptr_deref_1457_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1457_gather_scatter
    process(ptr_deref_1457_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1457_data_0;
      ov(7 downto 0) := iv;
      tmp44x_xi_1458 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1457_root_address_inst
    process(ptr_deref_1457_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1457_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1457_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1464_addr_0
    process(ptr_deref_1464_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1464_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1464_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1464_base_resize
    process(arrayidx48x_xi_1454) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx48x_xi_1454;
      ov := iv(2 downto 0);
      ptr_deref_1464_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1464_gather_scatter
    process(ptr_deref_1464_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1464_data_0;
      ov(7 downto 0) := iv;
      tmp49x_xi_1465 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1464_root_address_inst
    process(ptr_deref_1464_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1464_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1464_root_address <= ov(2 downto 0);
      --
    end process;
    if_stmt_1015_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1014;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1015_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1015_branch_req_0,
          ack0 => if_stmt_1015_branch_ack_0,
          ack1 => if_stmt_1015_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1177_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1176;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1177_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1177_branch_req_0,
          ack0 => if_stmt_1177_branch_ack_0,
          ack1 => if_stmt_1177_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1229_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1228;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1229_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1229_branch_req_0,
          ack0 => if_stmt_1229_branch_ack_0,
          ack1 => if_stmt_1229_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1383_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp53x_xi_1382;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1383_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1383_branch_req_0,
          ack0 => if_stmt_1383_branch_ack_0,
          ack1 => if_stmt_1383_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1480_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1479;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1480_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1480_branch_req_0,
          ack0 => if_stmt_1480_branch_ack_0,
          ack1 => if_stmt_1480_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1170_inst
    process(indvar_1049) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1049, type_cast_1169_wire_constant, tmp_var);
      indvarx_xnext_1171 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1400_inst
    process(and70_1222) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(and70_1222, type_cast_1399_wire_constant, tmp_var);
      tmpx_xopx_xi_1401 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1412_inst
    process(iNsTr_29_1407) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_29_1407, type_cast_1411_wire_constant, tmp_var);
      xx_xopx_xi_1413 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1447_inst
    process(tmp2_1436) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_1436, type_cast_1446_wire_constant, tmp_var);
      tmp3_1448 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1473_inst
    process(indvarx_xi_1423) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvarx_xi_1423, type_cast_1472_wire_constant, tmp_var);
      indvarx_xnextx_xi_1474 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1221_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(size_buffer, type_cast_1220_wire_constant, tmp_var);
      and70_1222 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1406_inst
    process(tmpx_xopx_xi_1401) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tmpx_xopx_xi_1401, type_cast_1405_wire_constant, tmp_var);
      iNsTr_29_1407 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1204_inst
    process(type_cast_1200_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1200_wire, type_cast_1203_wire_constant, tmp_var);
      ASHR_i64_i64_1204_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1381_inst
    process(conv74_1239) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv74_1239, type_cast_1380_wire_constant, tmp_var);
      cmp53x_xi_1382 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1175_inst
    process(indvarx_xnext_1171, umax4_1046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1171, umax4_1046, tmp_var);
      exitcond_1176 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1227_inst
    process(and70_1222) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and70_1222, type_cast_1226_wire_constant, tmp_var);
      tobool_1228 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1478_inst
    process(indvarx_xnextx_xi_1474, tmp58x_xi_1420) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnextx_xi_1474, tmp58x_xi_1420, tmp_var);
      exitcond1_1479 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1026_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_1025_wire_constant, tmp_var);
      shr_1027 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1076_inst
    process(tmp5_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_1067, type_cast_1075_wire_constant, tmp_var);
      shr11_1077 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1086_inst
    process(tmp5_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_1067, type_cast_1085_wire_constant, tmp_var);
      shr17_1087 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1096_inst
    process(tmp5_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_1067, type_cast_1095_wire_constant, tmp_var);
      shr23_1097 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1106_inst
    process(tmp5_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_1067, type_cast_1105_wire_constant, tmp_var);
      shr29_1107 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1116_inst
    process(tmp5_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_1067, type_cast_1115_wire_constant, tmp_var);
      shr35_1117 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1126_inst
    process(tmp5_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_1067, type_cast_1125_wire_constant, tmp_var);
      shr41_1127 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1136_inst
    process(tmp5_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_1067, type_cast_1135_wire_constant, tmp_var);
      shr47_1137 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1255_inst
    process(tmp1x_xi_1250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_1250, type_cast_1254_wire_constant, tmp_var);
      shrx_xi_1256 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1276_inst
    process(tmp1x_xi_1250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_1250, type_cast_1275_wire_constant, tmp_var);
      shr7x_xi_1277 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1297_inst
    process(tmp1x_xi_1250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_1250, type_cast_1296_wire_constant, tmp_var);
      shr13x_xi_1298 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1318_inst
    process(tmp1x_xi_1250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_1250, type_cast_1317_wire_constant, tmp_var);
      shr19x_xi_1319 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1339_inst
    process(tmp1x_xi_1250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_1250, type_cast_1338_wire_constant, tmp_var);
      shr25x_xi_1340 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1360_inst
    process(tmp1x_xi_1250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_1250, type_cast_1359_wire_constant, tmp_var);
      shr31x_xi_1361 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1435_inst
    process(indvarx_xi_1423) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvarx_xi_1423, type_cast_1434_wire_constant, tmp_var);
      tmp2_1436 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1195_inst
    process(umax_1190) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1190, type_cast_1194_wire_constant, tmp_var);
      tmp81_1196 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_1394_inst
    process(conv74_1239) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv74_1239, type_cast_1393_wire_constant, tmp_var);
      tmp55x_xi_1395 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1013_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_1012_wire_constant, tmp_var);
      cmp77_1014 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1032_inst
    process(shr_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_1027, type_cast_1031_wire_constant, tmp_var);
      tmp80_1033 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1038_inst
    process(shr_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_1027, type_cast_1037_wire_constant, tmp_var);
      tmp_1039 <= tmp_var; --
    end process;
    -- shared split operator group (32) : array_obj_ref_1061_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1060_scaled;
      array_obj_ref_1061_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1061_index_offset_req_0;
      array_obj_ref_1061_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1061_index_offset_req_1;
      array_obj_ref_1061_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : array_obj_ref_1244_index_offset 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1243_scaled;
      array_obj_ref_1244_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1244_index_offset_req_0;
      array_obj_ref_1244_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1244_index_offset_req_1;
      array_obj_ref_1244_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : array_obj_ref_1441_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_tmp2_1440_scaled;
      array_obj_ref_1441_final_offset <= data_out(2 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1441_index_offset_req_0;
      array_obj_ref_1441_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1441_index_offset_req_1;
      array_obj_ref_1441_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_1453_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_tmp3_1452_scaled;
      array_obj_ref_1453_final_offset <= data_out(2 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1453_index_offset_req_0;
      array_obj_ref_1453_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1453_index_offset_req_1;
      array_obj_ref_1453_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared load operator group (0) : ptr_deref_1066_load_0 ptr_deref_1249_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1066_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1249_load_0_req_0;
      ptr_deref_1066_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1249_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1066_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1249_load_0_req_1;
      ptr_deref_1066_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1249_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1066_word_address_0 & ptr_deref_1249_word_address_0;
      ptr_deref_1066_data_0 <= data_out(127 downto 64);
      ptr_deref_1249_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1457_load_0 ptr_deref_1464_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1457_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1464_load_0_req_0;
      ptr_deref_1457_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1464_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1457_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1464_load_0_req_1;
      ptr_deref_1457_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1464_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1457_word_address_0 & ptr_deref_1464_word_address_0;
      ptr_deref_1457_data_0 <= data_out(15 downto 8);
      ptr_deref_1464_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 3,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(2 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_1269_store_0 ptr_deref_1374_store_0 ptr_deref_1332_store_0 ptr_deref_1311_store_0 ptr_deref_1353_store_0 ptr_deref_1290_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(17 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_1269_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1374_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_1332_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1311_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1353_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1290_store_0_req_0;
      ptr_deref_1269_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1374_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_1332_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1311_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1353_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1290_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_1269_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1374_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_1332_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1311_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1353_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1290_store_0_req_1;
      ptr_deref_1269_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1374_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_1332_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1311_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1353_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1290_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1269_word_address_0 & ptr_deref_1374_word_address_0 & ptr_deref_1332_word_address_0 & ptr_deref_1311_word_address_0 & ptr_deref_1353_word_address_0 & ptr_deref_1290_word_address_0;
      data_in <= ptr_deref_1269_data_0 & ptr_deref_1374_data_0 & ptr_deref_1332_data_0 & ptr_deref_1311_data_0 & ptr_deref_1353_data_0 & ptr_deref_1290_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 3,
        data_width => 8,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(2 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 6,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1142_inst WPIPE_maxpool_output_pipe_1145_inst WPIPE_maxpool_output_pipe_1148_inst WPIPE_maxpool_output_pipe_1151_inst WPIPE_maxpool_output_pipe_1154_inst WPIPE_maxpool_output_pipe_1157_inst WPIPE_maxpool_output_pipe_1160_inst WPIPE_maxpool_output_pipe_1163_inst WPIPE_maxpool_output_pipe_1459_inst WPIPE_maxpool_output_pipe_1466_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal sample_req, sample_ack : BooleanArray( 9 downto 0);
      signal update_req, update_ack : BooleanArray( 9 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 9 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1142_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_1145_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1148_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1151_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1154_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1157_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1160_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1163_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1459_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1466_inst_req_0;
      WPIPE_maxpool_output_pipe_1142_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_1145_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_1148_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1151_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1154_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1157_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1160_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1163_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1459_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1466_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1142_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_1145_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1148_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1151_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1154_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1157_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1160_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1163_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1459_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1466_inst_req_1;
      WPIPE_maxpool_output_pipe_1142_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_1145_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_1148_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1151_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1154_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1157_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1160_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1163_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1459_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1466_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      data_in <= conv50_1141 & conv44_1131 & conv38_1121 & conv32_1111 & conv26_1101 & conv20_1091 & conv14_1081 & conv8_1071 & tmp44x_xi_1458 & tmp49x_xi_1465;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 10, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 3,
      data_width => 8,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 3,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendModule is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
    output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendModule;
architecture sendModule_arch of sendModule is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendModule_CP_8180_start: Boolean;
  signal sendModule_CP_8180_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal addr_of_3619_final_reg_req_1 : boolean;
  signal type_cast_3505_inst_req_0 : boolean;
  signal phi_stmt_3512_ack_0 : boolean;
  signal array_obj_ref_3628_index_offset_req_1 : boolean;
  signal addr_of_3629_final_reg_req_0 : boolean;
  signal addr_of_3629_final_reg_ack_1 : boolean;
  signal SUB_u16_u16_3531_inst_req_1 : boolean;
  signal addr_of_3629_final_reg_req_1 : boolean;
  signal addr_of_3629_final_reg_ack_0 : boolean;
  signal ptr_deref_3633_load_0_req_1 : boolean;
  signal ptr_deref_3633_load_0_ack_1 : boolean;
  signal addr_of_3619_final_reg_req_0 : boolean;
  signal phi_stmt_3507_req_0 : boolean;
  signal addr_of_3619_final_reg_ack_0 : boolean;
  signal array_obj_ref_3628_index_offset_ack_1 : boolean;
  signal SUB_u16_u16_3531_inst_ack_1 : boolean;
  signal type_cast_3505_inst_ack_1 : boolean;
  signal type_cast_3505_inst_req_1 : boolean;
  signal ptr_deref_3637_load_0_req_1 : boolean;
  signal ptr_deref_3637_load_0_ack_1 : boolean;
  signal array_obj_ref_3618_index_offset_ack_1 : boolean;
  signal array_obj_ref_3628_index_offset_ack_0 : boolean;
  signal ptr_deref_3637_load_0_req_0 : boolean;
  signal ptr_deref_3637_load_0_ack_0 : boolean;
  signal ptr_deref_3633_load_0_req_0 : boolean;
  signal ptr_deref_3633_load_0_ack_0 : boolean;
  signal array_obj_ref_3618_index_offset_req_1 : boolean;
  signal array_obj_ref_3628_index_offset_req_0 : boolean;
  signal n_row_3558_3521_buf_ack_1 : boolean;
  signal n_row_3558_3521_buf_req_1 : boolean;
  signal type_cast_3505_inst_ack_0 : boolean;
  signal phi_stmt_3517_ack_0 : boolean;
  signal array_obj_ref_3618_index_offset_ack_0 : boolean;
  signal addr_of_3619_final_reg_ack_1 : boolean;
  signal n_col_3547_3516_buf_ack_0 : boolean;
  signal phi_stmt_3517_req_0 : boolean;
  signal RPIPE_output_pipe_3481_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3481_inst_ack_0 : boolean;
  signal phi_stmt_3512_req_0 : boolean;
  signal RPIPE_output_pipe_3481_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3481_inst_ack_1 : boolean;
  signal type_cast_3569_inst_ack_0 : boolean;
  signal n_row_3558_3521_buf_ack_0 : boolean;
  signal RPIPE_output_pipe_3484_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3484_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3484_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3484_inst_ack_1 : boolean;
  signal array_obj_ref_3618_index_offset_req_0 : boolean;
  signal n_row_3558_3521_buf_req_0 : boolean;
  signal RPIPE_output_pipe_3487_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3487_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3487_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3487_inst_ack_1 : boolean;
  signal type_cast_3569_inst_req_0 : boolean;
  signal n_address2_3610_3506_buf_ack_1 : boolean;
  signal phi_stmt_3512_req_1 : boolean;
  signal do_while_stmt_3495_branch_req_0 : boolean;
  signal n_col_3547_3516_buf_req_0 : boolean;
  signal SUB_u16_u16_3531_inst_ack_0 : boolean;
  signal phi_stmt_3517_req_1 : boolean;
  signal type_cast_3569_inst_ack_1 : boolean;
  signal type_cast_3569_inst_req_1 : boolean;
  signal phi_stmt_3497_req_1 : boolean;
  signal phi_stmt_3497_req_0 : boolean;
  signal phi_stmt_3497_ack_0 : boolean;
  signal type_cast_3578_inst_ack_1 : boolean;
  signal n_col_3547_3516_buf_ack_1 : boolean;
  signal n_col_3547_3516_buf_req_1 : boolean;
  signal type_cast_3578_inst_req_1 : boolean;
  signal n_chl_3566_3511_buf_ack_1 : boolean;
  signal n_chl_3566_3511_buf_req_1 : boolean;
  signal n_chl_3566_3511_buf_ack_0 : boolean;
  signal n_chl_3566_3511_buf_req_0 : boolean;
  signal n_address1_3596_3501_buf_req_0 : boolean;
  signal phi_stmt_3507_ack_0 : boolean;
  signal n_address1_3596_3501_buf_ack_0 : boolean;
  signal n_address2_3610_3506_buf_req_1 : boolean;
  signal n_address1_3596_3501_buf_req_1 : boolean;
  signal n_address1_3596_3501_buf_ack_1 : boolean;
  signal type_cast_3578_inst_ack_0 : boolean;
  signal type_cast_3578_inst_req_0 : boolean;
  signal phi_stmt_3507_req_1 : boolean;
  signal SUB_u16_u16_3531_inst_req_0 : boolean;
  signal phi_stmt_3502_req_1 : boolean;
  signal n_address2_3610_3506_buf_ack_0 : boolean;
  signal phi_stmt_3502_req_0 : boolean;
  signal n_address2_3610_3506_buf_req_0 : boolean;
  signal phi_stmt_3502_ack_0 : boolean;
  signal RPIPE_output_pipe_3640_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3640_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3640_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3640_inst_ack_1 : boolean;
  signal RPIPE_output_pipe_3643_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3643_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3643_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3643_inst_ack_1 : boolean;
  signal slice_3647_inst_req_0 : boolean;
  signal slice_3647_inst_ack_0 : boolean;
  signal slice_3647_inst_req_1 : boolean;
  signal slice_3647_inst_ack_1 : boolean;
  signal slice_3651_inst_req_0 : boolean;
  signal slice_3651_inst_ack_0 : boolean;
  signal slice_3651_inst_req_1 : boolean;
  signal slice_3651_inst_ack_1 : boolean;
  signal slice_3655_inst_req_0 : boolean;
  signal slice_3655_inst_ack_0 : boolean;
  signal slice_3655_inst_req_1 : boolean;
  signal slice_3655_inst_ack_1 : boolean;
  signal slice_3659_inst_req_0 : boolean;
  signal slice_3659_inst_ack_0 : boolean;
  signal slice_3659_inst_req_1 : boolean;
  signal slice_3659_inst_ack_1 : boolean;
  signal slice_3663_inst_req_0 : boolean;
  signal slice_3663_inst_ack_0 : boolean;
  signal slice_3663_inst_req_1 : boolean;
  signal slice_3663_inst_ack_1 : boolean;
  signal slice_3667_inst_req_0 : boolean;
  signal slice_3667_inst_ack_0 : boolean;
  signal slice_3667_inst_req_1 : boolean;
  signal slice_3667_inst_ack_1 : boolean;
  signal slice_3671_inst_req_0 : boolean;
  signal slice_3671_inst_ack_0 : boolean;
  signal slice_3671_inst_req_1 : boolean;
  signal slice_3671_inst_ack_1 : boolean;
  signal slice_3675_inst_req_0 : boolean;
  signal slice_3675_inst_ack_0 : boolean;
  signal slice_3675_inst_req_1 : boolean;
  signal slice_3675_inst_ack_1 : boolean;
  signal W_output_data1_3560_delayed_14_0_3685_inst_req_0 : boolean;
  signal W_output_data1_3560_delayed_14_0_3685_inst_ack_0 : boolean;
  signal W_output_data1_3560_delayed_14_0_3685_inst_req_1 : boolean;
  signal W_output_data1_3560_delayed_14_0_3685_inst_ack_1 : boolean;
  signal EQ_u2_u1_3691_inst_req_0 : boolean;
  signal EQ_u2_u1_3691_inst_ack_0 : boolean;
  signal EQ_u2_u1_3691_inst_req_1 : boolean;
  signal EQ_u2_u1_3691_inst_ack_1 : boolean;
  signal EQ_u2_u1_3702_inst_req_0 : boolean;
  signal EQ_u2_u1_3702_inst_ack_0 : boolean;
  signal EQ_u2_u1_3702_inst_req_1 : boolean;
  signal EQ_u2_u1_3702_inst_ack_1 : boolean;
  signal W_output_data1_3568_delayed_14_0_3704_inst_req_0 : boolean;
  signal W_output_data1_3568_delayed_14_0_3704_inst_ack_0 : boolean;
  signal W_output_data1_3568_delayed_14_0_3704_inst_req_1 : boolean;
  signal W_output_data1_3568_delayed_14_0_3704_inst_ack_1 : boolean;
  signal EQ_u2_u1_3716_inst_req_0 : boolean;
  signal EQ_u2_u1_3716_inst_ack_0 : boolean;
  signal EQ_u2_u1_3716_inst_req_1 : boolean;
  signal EQ_u2_u1_3716_inst_ack_1 : boolean;
  signal W_output_data1_3576_delayed_14_0_3718_inst_req_0 : boolean;
  signal W_output_data1_3576_delayed_14_0_3718_inst_ack_0 : boolean;
  signal W_output_data1_3576_delayed_14_0_3718_inst_req_1 : boolean;
  signal W_output_data1_3576_delayed_14_0_3718_inst_ack_1 : boolean;
  signal EQ_u2_u1_3730_inst_req_0 : boolean;
  signal EQ_u2_u1_3730_inst_ack_0 : boolean;
  signal EQ_u2_u1_3730_inst_req_1 : boolean;
  signal EQ_u2_u1_3730_inst_ack_1 : boolean;
  signal W_output_data1_3584_delayed_14_0_3732_inst_req_0 : boolean;
  signal W_output_data1_3584_delayed_14_0_3732_inst_ack_0 : boolean;
  signal W_output_data1_3584_delayed_14_0_3732_inst_req_1 : boolean;
  signal W_output_data1_3584_delayed_14_0_3732_inst_ack_1 : boolean;
  signal EQ_u2_u1_3744_inst_req_0 : boolean;
  signal EQ_u2_u1_3744_inst_ack_0 : boolean;
  signal EQ_u2_u1_3744_inst_req_1 : boolean;
  signal EQ_u2_u1_3744_inst_ack_1 : boolean;
  signal W_output_data2_3592_delayed_14_0_3746_inst_req_0 : boolean;
  signal W_output_data2_3592_delayed_14_0_3746_inst_ack_0 : boolean;
  signal W_output_data2_3592_delayed_14_0_3746_inst_req_1 : boolean;
  signal W_output_data2_3592_delayed_14_0_3746_inst_ack_1 : boolean;
  signal EQ_u2_u1_3758_inst_req_0 : boolean;
  signal EQ_u2_u1_3758_inst_ack_0 : boolean;
  signal EQ_u2_u1_3758_inst_req_1 : boolean;
  signal EQ_u2_u1_3758_inst_ack_1 : boolean;
  signal W_output_data2_3600_delayed_14_0_3760_inst_req_0 : boolean;
  signal W_output_data2_3600_delayed_14_0_3760_inst_ack_0 : boolean;
  signal W_output_data2_3600_delayed_14_0_3760_inst_req_1 : boolean;
  signal W_output_data2_3600_delayed_14_0_3760_inst_ack_1 : boolean;
  signal EQ_u2_u1_3772_inst_req_0 : boolean;
  signal EQ_u2_u1_3772_inst_ack_0 : boolean;
  signal EQ_u2_u1_3772_inst_req_1 : boolean;
  signal EQ_u2_u1_3772_inst_ack_1 : boolean;
  signal W_output_data2_3608_delayed_14_0_3774_inst_req_0 : boolean;
  signal W_output_data2_3608_delayed_14_0_3774_inst_ack_0 : boolean;
  signal W_output_data2_3608_delayed_14_0_3774_inst_req_1 : boolean;
  signal W_output_data2_3608_delayed_14_0_3774_inst_ack_1 : boolean;
  signal EQ_u2_u1_3786_inst_req_0 : boolean;
  signal EQ_u2_u1_3786_inst_ack_0 : boolean;
  signal EQ_u2_u1_3786_inst_req_1 : boolean;
  signal EQ_u2_u1_3786_inst_ack_1 : boolean;
  signal W_output_data2_3616_delayed_14_0_3788_inst_req_0 : boolean;
  signal W_output_data2_3616_delayed_14_0_3788_inst_ack_0 : boolean;
  signal W_output_data2_3616_delayed_14_0_3788_inst_req_1 : boolean;
  signal W_output_data2_3616_delayed_14_0_3788_inst_ack_1 : boolean;
  signal W_fetch_addr1_3620_delayed_8_0_3797_inst_req_0 : boolean;
  signal W_fetch_addr1_3620_delayed_8_0_3797_inst_ack_0 : boolean;
  signal W_fetch_addr1_3620_delayed_8_0_3797_inst_req_1 : boolean;
  signal W_fetch_addr1_3620_delayed_8_0_3797_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3808_inst_req_0 : boolean;
  signal CONCAT_u32_u64_3808_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_3808_inst_req_1 : boolean;
  signal CONCAT_u32_u64_3808_inst_ack_1 : boolean;
  signal ptr_deref_3801_store_0_req_0 : boolean;
  signal ptr_deref_3801_store_0_ack_0 : boolean;
  signal ptr_deref_3801_store_0_req_1 : boolean;
  signal ptr_deref_3801_store_0_ack_1 : boolean;
  signal W_fetch_addr2_3630_delayed_8_0_3810_inst_req_0 : boolean;
  signal W_fetch_addr2_3630_delayed_8_0_3810_inst_ack_0 : boolean;
  signal W_fetch_addr2_3630_delayed_8_0_3810_inst_req_1 : boolean;
  signal W_fetch_addr2_3630_delayed_8_0_3810_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3821_inst_req_0 : boolean;
  signal CONCAT_u32_u64_3821_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_3821_inst_req_1 : boolean;
  signal CONCAT_u32_u64_3821_inst_ack_1 : boolean;
  signal ptr_deref_3814_store_0_req_0 : boolean;
  signal ptr_deref_3814_store_0_ack_0 : boolean;
  signal ptr_deref_3814_store_0_req_1 : boolean;
  signal ptr_deref_3814_store_0_ack_1 : boolean;
  signal SUB_u16_u16_3826_inst_req_0 : boolean;
  signal SUB_u16_u16_3826_inst_ack_0 : boolean;
  signal SUB_u16_u16_3826_inst_req_1 : boolean;
  signal SUB_u16_u16_3826_inst_ack_1 : boolean;
  signal do_while_stmt_3495_branch_ack_0 : boolean;
  signal do_while_stmt_3495_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3838_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3838_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_3838_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_3838_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendModule_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendModule_CP_8180_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendModule_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_8180_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendModule_CP_8180_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_8180_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendModule_CP_8180: Block -- control-path 
    signal sendModule_CP_8180_elements: BooleanArray(291 downto 0);
    -- 
  begin -- 
    sendModule_CP_8180_elements(0) <= sendModule_CP_8180_start;
    sendModule_CP_8180_symbol <= sendModule_CP_8180_elements(291);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3479/$entry
      -- CP-element group 0: 	 branch_block_stmt_3479/branch_block_stmt_3479__entry__
      -- CP-element group 0: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494__entry__
      -- CP-element group 0: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/$entry
      -- CP-element group 0: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_Sample/rr
      -- 
    rr_8204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(0), ack => RPIPE_output_pipe_3481_inst_req_0); -- 
    -- CP-element group 1:  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	289 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	290 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_3479/do_while_stmt_3495__exit__
      -- CP-element group 1: 	 branch_block_stmt_3479/assign_stmt_3840__entry__
      -- CP-element group 1: 	 branch_block_stmt_3479/assign_stmt_3840/$entry
      -- CP-element group 1: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_Sample/req
      -- 
    req_9281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(1), ack => WPIPE_input_done_pipe_3838_inst_req_0); -- 
    sendModule_CP_8180_elements(1) <= sendModule_CP_8180_elements(289);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_update_start_
      -- CP-element group 2: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_Update/cr
      -- 
    ra_8205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3481_inst_ack_0, ack => sendModule_CP_8180_elements(2)); -- 
    cr_8209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(2), ack => RPIPE_output_pipe_3481_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3481_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_Sample/rr
      -- 
    ca_8210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3481_inst_ack_1, ack => sendModule_CP_8180_elements(3)); -- 
    rr_8218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(3), ack => RPIPE_output_pipe_3484_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_update_start_
      -- CP-element group 4: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_Update/cr
      -- 
    ra_8219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3484_inst_ack_0, ack => sendModule_CP_8180_elements(4)); -- 
    cr_8223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(4), ack => RPIPE_output_pipe_3484_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3484_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_Sample/rr
      -- 
    ca_8224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3484_inst_ack_1, ack => sendModule_CP_8180_elements(5)); -- 
    rr_8232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(5), ack => RPIPE_output_pipe_3487_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_update_start_
      -- CP-element group 6: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_Update/cr
      -- 
    ra_8233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3487_inst_ack_0, ack => sendModule_CP_8180_elements(6)); -- 
    cr_8237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(6), ack => RPIPE_output_pipe_3487_inst_req_1); -- 
    -- CP-element group 7:  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494__exit__
      -- CP-element group 7: 	 branch_block_stmt_3479/do_while_stmt_3495__entry__
      -- CP-element group 7: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/$exit
      -- CP-element group 7: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_3479/assign_stmt_3482_to_assign_stmt_3494/RPIPE_output_pipe_3487_Update/ca
      -- 
    ca_8238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3487_inst_ack_1, ack => sendModule_CP_8180_elements(7)); -- 
    -- CP-element group 8:  transition  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_3479/do_while_stmt_3495/$entry
      -- CP-element group 8: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495__entry__
      -- 
    sendModule_CP_8180_elements(8) <= sendModule_CP_8180_elements(7);
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	289 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495__exit__
      -- 
    -- Element group sendModule_CP_8180_elements(9) is bound as output of CP function.
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3479/do_while_stmt_3495/loop_back
      -- 
    -- Element group sendModule_CP_8180_elements(10) is bound as output of CP function.
    -- CP-element group 11:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	287 
    -- CP-element group 11: 	288 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_3479/do_while_stmt_3495/condition_done
      -- CP-element group 11: 	 branch_block_stmt_3479/do_while_stmt_3495/loop_exit/$entry
      -- CP-element group 11: 	 branch_block_stmt_3479/do_while_stmt_3495/loop_taken/$entry
      -- 
    sendModule_CP_8180_elements(11) <= sendModule_CP_8180_elements(16);
    -- CP-element group 12:  branch  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	286 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_3479/do_while_stmt_3495/loop_body_done
      -- 
    sendModule_CP_8180_elements(12) <= sendModule_CP_8180_elements(286);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	65 
    -- CP-element group 13: 	84 
    -- CP-element group 13: 	103 
    -- CP-element group 13: 	25 
    -- CP-element group 13: 	44 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/back_edge_to_loop_body
      -- 
    sendModule_CP_8180_elements(13) <= sendModule_CP_8180_elements(10);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	67 
    -- CP-element group 14: 	86 
    -- CP-element group 14: 	105 
    -- CP-element group 14: 	27 
    -- CP-element group 14: 	46 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/first_time_through_loop_body
      -- 
    sendModule_CP_8180_elements(14) <= sendModule_CP_8180_elements(8);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	116 
    -- CP-element group 15: 	120 
    -- CP-element group 15: 	124 
    -- CP-element group 15: 	129 
    -- CP-element group 15: 	130 
    -- CP-element group 15: 	136 
    -- CP-element group 15: 	137 
    -- CP-element group 15: 	278 
    -- CP-element group 15: 	282 
    -- CP-element group 15: 	59 
    -- CP-element group 15: 	60 
    -- CP-element group 15: 	78 
    -- CP-element group 15: 	79 
    -- CP-element group 15: 	97 
    -- CP-element group 15: 	98 
    -- CP-element group 15: 	150 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	39 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/$entry
      -- CP-element group 15: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/loop_body_start
      -- 
    -- Element group sendModule_CP_8180_elements(15) is bound as output of CP function.
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	119 
    -- CP-element group 16: 	281 
    -- CP-element group 16: 	282 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/condition_evaluated
      -- 
    condition_evaluated_8253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_8253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(16), ack => do_while_stmt_3495_branch_req_0); -- 
    sendModule_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(20) & sendModule_CP_8180_elements(119) & sendModule_CP_8180_elements(281) & sendModule_CP_8180_elements(282);
      gj_sendModule_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	78 
    -- CP-element group 17: 	97 
    -- CP-element group 17: 	38 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	61 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	99 
    -- CP-element group 17: 	40 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/aggregated_phi_sample_req
      -- CP-element group 17: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_sample_start__ps
      -- 
    sendModule_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(21) & sendModule_CP_8180_elements(59) & sendModule_CP_8180_elements(78) & sendModule_CP_8180_elements(97) & sendModule_CP_8180_elements(38) & sendModule_CP_8180_elements(20);
      gj_sendModule_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	23 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	81 
    -- CP-element group 18: 	100 
    -- CP-element group 18: 	41 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	117 
    -- CP-element group 18: 	121 
    -- CP-element group 18: 	125 
    -- CP-element group 18: 	286 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	78 
    -- CP-element group 18: 	97 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/aggregated_phi_sample_ack
      -- CP-element group 18: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_sample_completed_
      -- 
    sendModule_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(23) & sendModule_CP_8180_elements(62) & sendModule_CP_8180_elements(81) & sendModule_CP_8180_elements(100) & sendModule_CP_8180_elements(41);
      gj_sendModule_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	60 
    -- CP-element group 19: 	79 
    -- CP-element group 19: 	98 
    -- CP-element group 19: 	39 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	63 
    -- CP-element group 19: 	82 
    -- CP-element group 19: 	101 
    -- CP-element group 19: 	42 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/aggregated_phi_update_req
      -- CP-element group 19: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_update_start__ps
      -- 
    sendModule_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(22) & sendModule_CP_8180_elements(60) & sendModule_CP_8180_elements(79) & sendModule_CP_8180_elements(98) & sendModule_CP_8180_elements(39);
      gj_sendModule_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	64 
    -- CP-element group 20: 	83 
    -- CP-element group 20: 	102 
    -- CP-element group 20: 	43 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/aggregated_phi_update_ack
      -- 
    sendModule_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(24) & sendModule_CP_8180_elements(64) & sendModule_CP_8180_elements(83) & sendModule_CP_8180_elements(102) & sendModule_CP_8180_elements(43);
      gj_sendModule_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	119 
    -- CP-element group 21: 	123 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_sample_start_
      -- 
    sendModule_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(18) & sendModule_CP_8180_elements(119) & sendModule_CP_8180_elements(123);
      gj_sendModule_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	196 
    -- CP-element group 22: 	200 
    -- CP-element group 22: 	208 
    -- CP-element group 22: 	216 
    -- CP-element group 22: 	131 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	19 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_update_start_
      -- 
    sendModule_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(196) & sendModule_CP_8180_elements(200) & sendModule_CP_8180_elements(208) & sendModule_CP_8180_elements(216) & sendModule_CP_8180_elements(131);
      gj_sendModule_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	18 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_sample_completed__ps
      -- 
    -- Element group sendModule_CP_8180_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	194 
    -- CP-element group 24: 	198 
    -- CP-element group 24: 	206 
    -- CP-element group 24: 	214 
    -- CP-element group 24: 	20 
    -- CP-element group 24: 	131 
    -- CP-element group 24:  members (15) 
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_scale_1/$entry
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_resize_1/index_resize_ack
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_resize_1/index_resize_req
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_scale_1/scale_rename_ack
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_resize_1/$exit
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_resize_1/$entry
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_Sample/req
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_computed_1
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_scale_1/scale_rename_req
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_scaled_1
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_resized_1
      -- CP-element group 24: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_index_scale_1/$exit
      -- 
    req_8555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(24), ack => array_obj_ref_3618_index_offset_req_0); -- 
    -- Element group sendModule_CP_8180_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	13 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_loopback_trigger
      -- 
    sendModule_CP_8180_elements(25) <= sendModule_CP_8180_elements(13);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_loopback_sample_req
      -- CP-element group 26: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_loopback_sample_req_ps
      -- 
    phi_stmt_3497_loopback_sample_req_8268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3497_loopback_sample_req_8268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(26), ack => phi_stmt_3497_req_1); -- 
    -- Element group sendModule_CP_8180_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	14 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_entry_trigger
      -- 
    sendModule_CP_8180_elements(27) <= sendModule_CP_8180_elements(14);
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_entry_sample_req
      -- CP-element group 28: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_entry_sample_req_ps
      -- 
    phi_stmt_3497_entry_sample_req_8271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3497_entry_sample_req_8271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(28), ack => phi_stmt_3497_req_0); -- 
    -- Element group sendModule_CP_8180_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_phi_mux_ack
      -- CP-element group 29: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3497_phi_mux_ack_ps
      -- 
    phi_stmt_3497_phi_mux_ack_8274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3497_ack_0, ack => sendModule_CP_8180_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3500_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3500_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3500_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3500_sample_completed_
      -- 
    -- Element group sendModule_CP_8180_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3500_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3500_update_start_
      -- 
    -- Element group sendModule_CP_8180_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3500_update_completed__ps
      -- 
    sendModule_CP_8180_elements(32) <= sendModule_CP_8180_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3500_update_completed_
      -- 
    -- Element group sendModule_CP_8180_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => sendModule_CP_8180_elements(31), ack => sendModule_CP_8180_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_Sample/req
      -- 
    req_8295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(34), ack => n_address1_3596_3501_buf_req_0); -- 
    -- Element group sendModule_CP_8180_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_update_start_
      -- CP-element group 35: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_Update/req
      -- 
    req_8300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(35), ack => n_address1_3596_3501_buf_req_1); -- 
    -- Element group sendModule_CP_8180_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_Sample/ack
      -- 
    ack_8296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_3596_3501_buf_ack_0, ack => sendModule_CP_8180_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address1_3501_Update/ack
      -- 
    ack_8301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_3596_3501_buf_ack_1, ack => sendModule_CP_8180_elements(37)); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	18 
    -- CP-element group 38: 	119 
    -- CP-element group 38: 	127 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	17 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_sample_start_
      -- 
    sendModule_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(18) & sendModule_CP_8180_elements(119) & sendModule_CP_8180_elements(127);
      gj_sendModule_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	15 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	248 
    -- CP-element group 39: 	224 
    -- CP-element group 39: 	232 
    -- CP-element group 39: 	240 
    -- CP-element group 39: 	138 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	19 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_update_start_
      -- 
    sendModule_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(248) & sendModule_CP_8180_elements(224) & sendModule_CP_8180_elements(232) & sendModule_CP_8180_elements(240) & sendModule_CP_8180_elements(138);
      gj_sendModule_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	17 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_sample_start__ps
      -- 
    sendModule_CP_8180_elements(40) <= sendModule_CP_8180_elements(17);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	18 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_sample_completed__ps
      -- 
    -- Element group sendModule_CP_8180_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_update_start__ps
      -- 
    sendModule_CP_8180_elements(42) <= sendModule_CP_8180_elements(19);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	246 
    -- CP-element group 43: 	222 
    -- CP-element group 43: 	230 
    -- CP-element group 43: 	238 
    -- CP-element group 43: 	20 
    -- CP-element group 43: 	138 
    -- CP-element group 43:  members (15) 
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_scale_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_Sample/req
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_update_completed__ps
      -- 
    req_8601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(43), ack => array_obj_ref_3628_index_offset_req_0); -- 
    -- Element group sendModule_CP_8180_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	13 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_loopback_trigger
      -- 
    sendModule_CP_8180_elements(44) <= sendModule_CP_8180_elements(13);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_loopback_sample_req_ps
      -- 
    phi_stmt_3502_loopback_sample_req_8312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3502_loopback_sample_req_8312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(45), ack => phi_stmt_3502_req_1); -- 
    -- Element group sendModule_CP_8180_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	14 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_entry_trigger
      -- 
    sendModule_CP_8180_elements(46) <= sendModule_CP_8180_elements(14);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_entry_sample_req
      -- CP-element group 47: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_entry_sample_req_ps
      -- 
    phi_stmt_3502_entry_sample_req_8315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3502_entry_sample_req_8315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(47), ack => phi_stmt_3502_req_0); -- 
    -- Element group sendModule_CP_8180_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_phi_mux_ack
      -- CP-element group 48: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3502_phi_mux_ack_ps
      -- 
    phi_stmt_3502_phi_mux_ack_8318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3502_ack_0, ack => sendModule_CP_8180_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_sample_start__ps
      -- 
    -- Element group sendModule_CP_8180_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_update_start__ps
      -- 
    -- Element group sendModule_CP_8180_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_sample_start_
      -- 
    rr_8331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(51), ack => type_cast_3505_inst_req_0); -- 
    sendModule_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(49) & sendModule_CP_8180_elements(53);
      gj_sendModule_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_update_start_
      -- 
    cr_8336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(52), ack => type_cast_3505_inst_req_1); -- 
    sendModule_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(50) & sendModule_CP_8180_elements(54);
      gj_sendModule_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_sample_completed__ps
      -- 
    ra_8332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3505_inst_ack_0, ack => sendModule_CP_8180_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3505_update_completed__ps
      -- 
    ca_8337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3505_inst_ack_1, ack => sendModule_CP_8180_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_Sample/req
      -- 
    req_8349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(55), ack => n_address2_3610_3506_buf_req_0); -- 
    -- Element group sendModule_CP_8180_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_update_start_
      -- CP-element group 56: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_update_start__ps
      -- CP-element group 56: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_Update/req
      -- CP-element group 56: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_Update/$entry
      -- 
    req_8354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(56), ack => n_address2_3610_3506_buf_req_1); -- 
    -- Element group sendModule_CP_8180_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_Sample/ack
      -- 
    ack_8350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_3610_3506_buf_ack_0, ack => sendModule_CP_8180_elements(57)); -- 
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_address2_3506_Update/$exit
      -- 
    ack_8355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_3610_3506_buf_ack_1, ack => sendModule_CP_8180_elements(58)); -- 
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	15 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	119 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_sample_start_
      -- 
    sendModule_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(18) & sendModule_CP_8180_elements(119);
      gj_sendModule_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	15 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	64 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	19 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_update_start_
      -- 
    sendModule_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(64);
      gj_sendModule_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	17 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_sample_start__ps
      -- 
    sendModule_CP_8180_elements(61) <= sendModule_CP_8180_elements(17);
    -- CP-element group 62:  join  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	18 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_sample_completed__ps
      -- 
    -- Element group sendModule_CP_8180_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_update_start__ps
      -- 
    sendModule_CP_8180_elements(63) <= sendModule_CP_8180_elements(19);
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	20 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	60 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_update_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_update_completed_
      -- 
    -- Element group sendModule_CP_8180_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	13 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_loopback_trigger
      -- 
    sendModule_CP_8180_elements(65) <= sendModule_CP_8180_elements(13);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_loopback_sample_req_ps
      -- CP-element group 66: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_loopback_sample_req
      -- 
    phi_stmt_3507_loopback_sample_req_8366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3507_loopback_sample_req_8366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(66), ack => phi_stmt_3507_req_1); -- 
    -- Element group sendModule_CP_8180_elements(66) is bound as output of CP function.
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_entry_trigger
      -- 
    sendModule_CP_8180_elements(67) <= sendModule_CP_8180_elements(14);
    -- CP-element group 68:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_entry_sample_req
      -- CP-element group 68: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_entry_sample_req_ps
      -- 
    phi_stmt_3507_entry_sample_req_8369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3507_entry_sample_req_8369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(68), ack => phi_stmt_3507_req_0); -- 
    -- Element group sendModule_CP_8180_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_phi_mux_ack_ps
      -- CP-element group 69: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3507_phi_mux_ack
      -- 
    phi_stmt_3507_phi_mux_ack_8372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3507_ack_0, ack => sendModule_CP_8180_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3510_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3510_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3510_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3510_sample_start__ps
      -- 
    -- Element group sendModule_CP_8180_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3510_update_start_
      -- CP-element group 71: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3510_update_start__ps
      -- 
    -- Element group sendModule_CP_8180_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3510_update_completed__ps
      -- 
    sendModule_CP_8180_elements(72) <= sendModule_CP_8180_elements(73);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	72 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3510_update_completed_
      -- 
    -- Element group sendModule_CP_8180_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => sendModule_CP_8180_elements(71), ack => sendModule_CP_8180_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_sample_start__ps
      -- CP-element group 74: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_Sample/req
      -- 
    req_8393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(74), ack => n_chl_3566_3511_buf_req_0); -- 
    -- Element group sendModule_CP_8180_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_update_start_
      -- CP-element group 75: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_update_start__ps
      -- CP-element group 75: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_Update/req
      -- CP-element group 75: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_Update/$entry
      -- 
    req_8398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(75), ack => n_chl_3566_3511_buf_req_1); -- 
    -- Element group sendModule_CP_8180_elements(75) is bound as output of CP function.
    -- CP-element group 76:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_Sample/ack
      -- CP-element group 76: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_Sample/$exit
      -- 
    ack_8394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3566_3511_buf_ack_0, ack => sendModule_CP_8180_elements(76)); -- 
    -- CP-element group 77:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_Update/ack
      -- CP-element group 77: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_chl_3511_Update/$exit
      -- 
    ack_8399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3566_3511_buf_ack_1, ack => sendModule_CP_8180_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	15 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	18 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	17 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_sample_start_
      -- 
    sendModule_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(18);
      gj_sendModule_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	15 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	19 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_update_start_
      -- 
    sendModule_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(83);
      gj_sendModule_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_sample_start__ps
      -- 
    sendModule_CP_8180_elements(80) <= sendModule_CP_8180_elements(17);
    -- CP-element group 81:  join  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	18 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_sample_completed__ps
      -- 
    -- Element group sendModule_CP_8180_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	19 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_update_start__ps
      -- 
    sendModule_CP_8180_elements(82) <= sendModule_CP_8180_elements(19);
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	20 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_update_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_update_completed_
      -- 
    -- Element group sendModule_CP_8180_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	13 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_loopback_trigger
      -- 
    sendModule_CP_8180_elements(84) <= sendModule_CP_8180_elements(13);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_loopback_sample_req_ps
      -- CP-element group 85: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_loopback_sample_req
      -- 
    phi_stmt_3512_loopback_sample_req_8410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3512_loopback_sample_req_8410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(85), ack => phi_stmt_3512_req_1); -- 
    -- Element group sendModule_CP_8180_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	14 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_entry_trigger
      -- 
    sendModule_CP_8180_elements(86) <= sendModule_CP_8180_elements(14);
    -- CP-element group 87:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_entry_sample_req_ps
      -- CP-element group 87: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_entry_sample_req
      -- 
    phi_stmt_3512_entry_sample_req_8413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3512_entry_sample_req_8413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(87), ack => phi_stmt_3512_req_0); -- 
    -- Element group sendModule_CP_8180_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_phi_mux_ack
      -- CP-element group 88: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3512_phi_mux_ack_ps
      -- 
    phi_stmt_3512_phi_mux_ack_8416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3512_ack_0, ack => sendModule_CP_8180_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3515_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3515_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3515_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3515_sample_start__ps
      -- 
    -- Element group sendModule_CP_8180_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3515_update_start_
      -- CP-element group 90: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3515_update_start__ps
      -- 
    -- Element group sendModule_CP_8180_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3515_update_completed__ps
      -- 
    sendModule_CP_8180_elements(91) <= sendModule_CP_8180_elements(92);
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3515_update_completed_
      -- 
    -- Element group sendModule_CP_8180_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => sendModule_CP_8180_elements(90), ack => sendModule_CP_8180_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_sample_start__ps
      -- CP-element group 93: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_Sample/req
      -- CP-element group 93: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_Sample/$entry
      -- 
    req_8437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(93), ack => n_col_3547_3516_buf_req_0); -- 
    -- Element group sendModule_CP_8180_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_update_start__ps
      -- CP-element group 94: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_Update/req
      -- CP-element group 94: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_update_start_
      -- 
    req_8442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(94), ack => n_col_3547_3516_buf_req_1); -- 
    -- Element group sendModule_CP_8180_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_Sample/ack
      -- CP-element group 95: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_sample_completed_
      -- 
    ack_8438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3547_3516_buf_ack_0, ack => sendModule_CP_8180_elements(95)); -- 
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_Update/ack
      -- CP-element group 96: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_col_3516_Update/$exit
      -- 
    ack_8443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3547_3516_buf_ack_1, ack => sendModule_CP_8180_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	15 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	18 
    -- CP-element group 97: 	119 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	17 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_sample_start_
      -- 
    sendModule_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(18) & sendModule_CP_8180_elements(119);
      gj_sendModule_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	15 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	19 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_update_start_
      -- 
    sendModule_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(102);
      gj_sendModule_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	17 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_sample_start__ps
      -- 
    sendModule_CP_8180_elements(99) <= sendModule_CP_8180_elements(17);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	18 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_sample_completed__ps
      -- 
    -- Element group sendModule_CP_8180_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	19 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_update_start__ps
      -- 
    sendModule_CP_8180_elements(101) <= sendModule_CP_8180_elements(19);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	20 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_update_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_update_completed_
      -- 
    -- Element group sendModule_CP_8180_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	13 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_loopback_trigger
      -- 
    sendModule_CP_8180_elements(103) <= sendModule_CP_8180_elements(13);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_loopback_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_loopback_sample_req
      -- 
    phi_stmt_3517_loopback_sample_req_8454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3517_loopback_sample_req_8454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(104), ack => phi_stmt_3517_req_1); -- 
    -- Element group sendModule_CP_8180_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	14 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_entry_trigger
      -- 
    sendModule_CP_8180_elements(105) <= sendModule_CP_8180_elements(14);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_entry_sample_req_ps
      -- CP-element group 106: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_entry_sample_req
      -- 
    phi_stmt_3517_entry_sample_req_8457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3517_entry_sample_req_8457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(106), ack => phi_stmt_3517_req_0); -- 
    -- Element group sendModule_CP_8180_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_phi_mux_ack_ps
      -- CP-element group 107: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/phi_stmt_3517_phi_mux_ack
      -- 
    phi_stmt_3517_phi_mux_ack_8460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3517_ack_0, ack => sendModule_CP_8180_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3520_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3520_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3520_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3520_sample_start__ps
      -- 
    -- Element group sendModule_CP_8180_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3520_update_start_
      -- CP-element group 109: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3520_update_start__ps
      -- 
    -- Element group sendModule_CP_8180_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3520_update_completed__ps
      -- 
    sendModule_CP_8180_elements(110) <= sendModule_CP_8180_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3520_update_completed_
      -- 
    -- Element group sendModule_CP_8180_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => sendModule_CP_8180_elements(109), ack => sendModule_CP_8180_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_Sample/req
      -- CP-element group 112: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_sample_start__ps
      -- 
    req_8481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(112), ack => n_row_3558_3521_buf_req_0); -- 
    -- Element group sendModule_CP_8180_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_Update/req
      -- CP-element group 113: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_update_start_
      -- CP-element group 113: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_update_start__ps
      -- 
    req_8486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(113), ack => n_row_3558_3521_buf_req_1); -- 
    -- Element group sendModule_CP_8180_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_sample_completed__ps
      -- 
    ack_8482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3558_3521_buf_ack_0, ack => sendModule_CP_8180_elements(114)); -- 
    -- CP-element group 115:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_Update/ack
      -- CP-element group 115: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/R_n_row_3521_update_completed__ps
      -- 
    ack_8487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3558_3521_buf_ack_1, ack => sendModule_CP_8180_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	15 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_Sample/$entry
      -- 
    rr_8496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(116), ack => SUB_u16_u16_3531_inst_req_0); -- 
    sendModule_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(118);
      gj_sendModule_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	18 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_update_start_
      -- CP-element group 117: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_Update/cr
      -- CP-element group 117: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_Update/$entry
      -- 
    cr_8501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(117), ack => SUB_u16_u16_3531_inst_req_1); -- 
    sendModule_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(18) & sendModule_CP_8180_elements(119);
      gj_sendModule_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_Sample/$exit
      -- 
    ra_8497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3531_inst_ack_0, ack => sendModule_CP_8180_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	16 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	21 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	59 
    -- CP-element group 119: 	97 
    -- CP-element group 119: 	38 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3531_Update/$exit
      -- 
    ca_8502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3531_inst_ack_1, ack => sendModule_CP_8180_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	15 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_Sample/$entry
      -- 
    rr_8510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(120), ack => type_cast_3569_inst_req_0); -- 
    sendModule_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(122);
      gj_sendModule_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	18 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_update_start_
      -- CP-element group 121: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_Update/cr
      -- 
    cr_8515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(121), ack => type_cast_3569_inst_req_1); -- 
    sendModule_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(18) & sendModule_CP_8180_elements(123);
      gj_sendModule_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_Sample/$exit
      -- 
    ra_8511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3569_inst_ack_0, ack => sendModule_CP_8180_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	286 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	21 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3569_Update/ca
      -- 
    ca_8516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3569_inst_ack_1, ack => sendModule_CP_8180_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	15 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_Sample/rr
      -- CP-element group 124: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_Sample/$entry
      -- 
    rr_8524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(124), ack => type_cast_3578_inst_req_0); -- 
    sendModule_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(126);
      gj_sendModule_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	18 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_update_start_
      -- CP-element group 125: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_Update/cr
      -- CP-element group 125: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_Update/$entry
      -- 
    cr_8529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(125), ack => type_cast_3578_inst_req_1); -- 
    sendModule_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(18) & sendModule_CP_8180_elements(127);
      gj_sendModule_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_Sample/ra
      -- CP-element group 126: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_Sample/$exit
      -- 
    ra_8525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3578_inst_ack_0, ack => sendModule_CP_8180_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	286 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	38 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/type_cast_3578_update_completed_
      -- 
    ca_8530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3578_inst_ack_1, ack => sendModule_CP_8180_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	132 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	133 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_request/req
      -- CP-element group 128: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_request/$entry
      -- CP-element group 128: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_sample_start_
      -- 
    req_8570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(128), ack => addr_of_3619_final_reg_req_0); -- 
    sendModule_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(132) & sendModule_CP_8180_elements(133);
      gj_sendModule_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	15 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	256 
    -- CP-element group 129: 	144 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	134 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_complete/req
      -- CP-element group 129: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_complete/$entry
      -- CP-element group 129: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_update_start_
      -- 
    req_8575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(129), ack => addr_of_3619_final_reg_req_1); -- 
    sendModule_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(256) & sendModule_CP_8180_elements(144);
      gj_sendModule_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	15 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	133 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_Update/req
      -- CP-element group 130: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_update_start
      -- CP-element group 130: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_Update/$entry
      -- 
    req_8560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(130), ack => array_obj_ref_3618_index_offset_req_1); -- 
    sendModule_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(133);
      gj_sendModule_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	24 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	286 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	22 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_sample_complete
      -- CP-element group 131: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_Sample/ack
      -- 
    ack_8556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3618_index_offset_ack_0, ack => sendModule_CP_8180_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	128 
    -- CP-element group 132:  members (8) 
      -- CP-element group 132: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_root_address_calculated
      -- CP-element group 132: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_Update/ack
      -- CP-element group 132: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_final_index_sum_regn_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_base_plus_offset/sum_rename_ack
      -- CP-element group 132: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_base_plus_offset/sum_rename_req
      -- CP-element group 132: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_base_plus_offset/$exit
      -- CP-element group 132: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_base_plus_offset/$entry
      -- CP-element group 132: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3618_offset_calculated
      -- 
    ack_8561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3618_index_offset_ack_1, ack => sendModule_CP_8180_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	130 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_request/ack
      -- CP-element group 133: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_request/$exit
      -- CP-element group 133: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_sample_completed_
      -- 
    ack_8571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3619_final_reg_ack_0, ack => sendModule_CP_8180_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	129 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	254 
    -- CP-element group 134: 	142 
    -- CP-element group 134:  members (19) 
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_plus_offset/$entry
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_addr_resize/$entry
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_word_addrgen/$exit
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_root_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_plus_offset/sum_rename_req
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_complete/$exit
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_word_addrgen/root_register_ack
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_word_addrgen/$entry
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_plus_offset/sum_rename_ack
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_addr_resize/base_resize_req
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_addr_resize/base_resize_ack
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_word_addrgen/root_register_req
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_address_resized
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_word_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_addr_resize/$exit
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_complete/ack
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3619_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_base_plus_offset/$exit
      -- 
    ack_8576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3619_final_reg_ack_1, ack => sendModule_CP_8180_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	139 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	140 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	140 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_request/$entry
      -- CP-element group 135: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_request/req
      -- 
    req_8616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(135), ack => addr_of_3629_final_reg_req_0); -- 
    sendModule_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(139) & sendModule_CP_8180_elements(140);
      gj_sendModule_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	15 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	268 
    -- CP-element group 136: 	148 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	141 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_update_start_
      -- CP-element group 136: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_complete/req
      -- CP-element group 136: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_complete/$entry
      -- 
    req_8621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(136), ack => addr_of_3629_final_reg_req_1); -- 
    sendModule_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(268) & sendModule_CP_8180_elements(148);
      gj_sendModule_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	15 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	140 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_Update/req
      -- CP-element group 137: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_update_start
      -- CP-element group 137: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_Update/$entry
      -- 
    req_8606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(137), ack => array_obj_ref_3628_index_offset_req_1); -- 
    sendModule_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(140);
      gj_sendModule_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	43 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	286 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	39 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_sample_complete
      -- CP-element group 138: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_Sample/ack
      -- CP-element group 138: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_Sample/$exit
      -- 
    ack_8602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3628_index_offset_ack_0, ack => sendModule_CP_8180_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	135 
    -- CP-element group 139:  members (8) 
      -- CP-element group 139: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_Update/ack
      -- CP-element group 139: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_base_plus_offset/$entry
      -- CP-element group 139: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_base_plus_offset/$exit
      -- CP-element group 139: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_final_index_sum_regn_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_offset_calculated
      -- CP-element group 139: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_base_plus_offset/sum_rename_ack
      -- CP-element group 139: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/array_obj_ref_3628_base_plus_offset/sum_rename_req
      -- 
    ack_8607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3628_index_offset_ack_1, ack => sendModule_CP_8180_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	135 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	135 
    -- CP-element group 140: 	137 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_request/$exit
      -- CP-element group 140: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_request/ack
      -- 
    ack_8617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3629_final_reg_ack_0, ack => sendModule_CP_8180_elements(140)); -- 
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	136 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	266 
    -- CP-element group 141: 	146 
    -- CP-element group 141:  members (19) 
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_complete/ack
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_complete/$exit
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_address_resized
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/addr_of_3629_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_word_addrgen/root_register_req
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_word_addrgen/root_register_ack
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_addr_resize/base_resize_req
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_addr_resize/base_resize_ack
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_addr_resize/$entry
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_addr_resize/$exit
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_word_addrgen/$entry
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_word_addrgen/$exit
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_base_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_word_address_calculated
      -- 
    ack_8622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3629_final_reg_ack_1, ack => sendModule_CP_8180_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	134 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	276 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (5) 
      -- CP-element group 142: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Sample/word_access_start/$entry
      -- CP-element group 142: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Sample/word_access_start/word_0/rr
      -- CP-element group 142: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Sample/word_access_start/word_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Sample/$entry
      -- 
    rr_8655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(142), ack => ptr_deref_3633_load_0_req_0); -- 
    sendModule_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(134) & sendModule_CP_8180_elements(276);
      gj_sendModule_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	160 
    -- CP-element group 143: 	164 
    -- CP-element group 143: 	168 
    -- CP-element group 143: 	172 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/word_access_complete/word_0/cr
      -- CP-element group 143: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/word_access_complete/$entry
      -- CP-element group 143: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_update_start_
      -- CP-element group 143: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/word_access_complete/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/$entry
      -- 
    cr_8666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(143), ack => ptr_deref_3633_load_0_req_1); -- 
    sendModule_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(160) & sendModule_CP_8180_elements(164) & sendModule_CP_8180_elements(168) & sendModule_CP_8180_elements(172);
      gj_sendModule_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	283 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	129 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Sample/word_access_start/word_0/ra
      -- CP-element group 144: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Sample/word_access_start/word_0/$exit
      -- 
    ra_8656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3633_load_0_ack_0, ack => sendModule_CP_8180_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	158 
    -- CP-element group 145: 	162 
    -- CP-element group 145: 	166 
    -- CP-element group 145: 	170 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/word_access_complete/word_0/ca
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/ptr_deref_3633_Merge/$entry
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/ptr_deref_3633_Merge/$exit
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/ptr_deref_3633_Merge/merge_req
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/ptr_deref_3633_Merge/merge_ack
      -- CP-element group 145: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_Update/$exit
      -- 
    ca_8667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3633_load_0_ack_1, ack => sendModule_CP_8180_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	141 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	276 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Sample/word_access_start/$entry
      -- CP-element group 146: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Sample/word_access_start/word_0/$entry
      -- CP-element group 146: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Sample/word_access_start/word_0/rr
      -- CP-element group 146: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Sample/$entry
      -- 
    rr_8705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(146), ack => ptr_deref_3637_load_0_req_0); -- 
    sendModule_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(141) & sendModule_CP_8180_elements(276);
      gj_sendModule_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	180 
    -- CP-element group 147: 	184 
    -- CP-element group 147: 	188 
    -- CP-element group 147: 	176 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_update_start_
      -- CP-element group 147: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/word_access_complete/word_0/cr
      -- CP-element group 147: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/word_access_complete/$entry
      -- CP-element group 147: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/word_access_complete/word_0/$entry
      -- 
    cr_8716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(147), ack => ptr_deref_3637_load_0_req_1); -- 
    sendModule_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(180) & sendModule_CP_8180_elements(184) & sendModule_CP_8180_elements(188) & sendModule_CP_8180_elements(176);
      gj_sendModule_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	284 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	136 
    -- CP-element group 148:  members (5) 
      -- CP-element group 148: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Sample/word_access_start/$exit
      -- CP-element group 148: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Sample/word_access_start/word_0/$exit
      -- CP-element group 148: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Sample/word_access_start/word_0/ra
      -- CP-element group 148: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Sample/$exit
      -- 
    ra_8706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3637_load_0_ack_0, ack => sendModule_CP_8180_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	182 
    -- CP-element group 149: 	186 
    -- CP-element group 149: 	174 
    -- CP-element group 149: 	178 
    -- CP-element group 149:  members (9) 
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/word_access_complete/word_0/$exit
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/word_access_complete/word_0/ca
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/ptr_deref_3637_Merge/$entry
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/word_access_complete/$exit
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/ptr_deref_3637_Merge/$exit
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/ptr_deref_3637_Merge/merge_req
      -- CP-element group 149: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_Update/ptr_deref_3637_Merge/merge_ack
      -- 
    ca_8717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3637_load_0_ack_1, ack => sendModule_CP_8180_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	15 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_Sample/rr
      -- 
    rr_8730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(150), ack => RPIPE_output_pipe_3640_inst_req_0); -- 
    sendModule_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(153);
      gj_sendModule_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	192 
    -- CP-element group 151: 	204 
    -- CP-element group 151: 	212 
    -- CP-element group 151: 	220 
    -- CP-element group 151: 	157 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_update_start_
      -- CP-element group 151: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_Update/cr
      -- 
    cr_8735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(151), ack => RPIPE_output_pipe_3640_inst_req_1); -- 
    sendModule_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(152) & sendModule_CP_8180_elements(192) & sendModule_CP_8180_elements(204) & sendModule_CP_8180_elements(212) & sendModule_CP_8180_elements(220) & sendModule_CP_8180_elements(157);
      gj_sendModule_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	151 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_Sample/ra
      -- 
    ra_8731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3640_inst_ack_0, ack => sendModule_CP_8180_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	190 
    -- CP-element group 153: 	202 
    -- CP-element group 153: 	210 
    -- CP-element group 153: 	218 
    -- CP-element group 153: 	154 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3640_Update/ca
      -- 
    ca_8736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3640_inst_ack_1, ack => sendModule_CP_8180_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	157 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_Sample/rr
      -- 
    rr_8744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(154), ack => RPIPE_output_pipe_3643_inst_req_0); -- 
    sendModule_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(153) & sendModule_CP_8180_elements(157);
      gj_sendModule_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	244 
    -- CP-element group 155: 	252 
    -- CP-element group 155: 	228 
    -- CP-element group 155: 	236 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_update_start_
      -- CP-element group 155: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_Update/cr
      -- 
    cr_8749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(155), ack => RPIPE_output_pipe_3643_inst_req_1); -- 
    sendModule_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(156) & sendModule_CP_8180_elements(244) & sendModule_CP_8180_elements(252) & sendModule_CP_8180_elements(228) & sendModule_CP_8180_elements(236);
      gj_sendModule_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	155 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_Sample/ra
      -- 
    ra_8745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3643_inst_ack_0, ack => sendModule_CP_8180_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	242 
    -- CP-element group 157: 	250 
    -- CP-element group 157: 	226 
    -- CP-element group 157: 	234 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	151 
    -- CP-element group 157: 	154 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/RPIPE_output_pipe_3643_Update/ca
      -- 
    ca_8750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3643_inst_ack_1, ack => sendModule_CP_8180_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	145 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_Sample/rr
      -- 
    rr_8758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(158), ack => slice_3647_inst_req_0); -- 
    sendModule_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(145) & sendModule_CP_8180_elements(160);
      gj_sendModule_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	260 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_update_start_
      -- CP-element group 159: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_Update/cr
      -- 
    cr_8763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(159), ack => slice_3647_inst_req_1); -- 
    sendModule_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	143 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_Sample/ra
      -- 
    ra_8759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3647_inst_ack_0, ack => sendModule_CP_8180_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	258 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3647_Update/ca
      -- 
    ca_8764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3647_inst_ack_1, ack => sendModule_CP_8180_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	145 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_Sample/rr
      -- 
    rr_8772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(162), ack => slice_3651_inst_req_0); -- 
    sendModule_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(145) & sendModule_CP_8180_elements(164);
      gj_sendModule_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	260 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_Update/cr
      -- 
    cr_8777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(163), ack => slice_3651_inst_req_1); -- 
    sendModule_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	143 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_Sample/ra
      -- 
    ra_8773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3651_inst_ack_0, ack => sendModule_CP_8180_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	258 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3651_Update/ca
      -- 
    ca_8778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3651_inst_ack_1, ack => sendModule_CP_8180_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	145 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_Sample/rr
      -- 
    rr_8786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(166), ack => slice_3655_inst_req_0); -- 
    sendModule_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(145) & sendModule_CP_8180_elements(168);
      gj_sendModule_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	260 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_update_start_
      -- CP-element group 167: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_Update/cr
      -- 
    cr_8791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(167), ack => slice_3655_inst_req_1); -- 
    sendModule_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	143 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_Sample/ra
      -- 
    ra_8787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3655_inst_ack_0, ack => sendModule_CP_8180_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	258 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3655_Update/ca
      -- 
    ca_8792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3655_inst_ack_1, ack => sendModule_CP_8180_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	145 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_Sample/rr
      -- 
    rr_8800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(170), ack => slice_3659_inst_req_0); -- 
    sendModule_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(145) & sendModule_CP_8180_elements(172);
      gj_sendModule_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	260 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_update_start_
      -- CP-element group 171: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_Update/cr
      -- 
    cr_8805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(171), ack => slice_3659_inst_req_1); -- 
    sendModule_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	143 
    -- CP-element group 172: 	170 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_Sample/ra
      -- 
    ra_8801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3659_inst_ack_0, ack => sendModule_CP_8180_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	258 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3659_Update/ca
      -- 
    ca_8806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3659_inst_ack_1, ack => sendModule_CP_8180_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	149 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_Sample/rr
      -- 
    rr_8814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(174), ack => slice_3663_inst_req_0); -- 
    sendModule_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(149) & sendModule_CP_8180_elements(176);
      gj_sendModule_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	272 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_update_start_
      -- CP-element group 175: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_Update/cr
      -- 
    cr_8819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(175), ack => slice_3663_inst_req_1); -- 
    sendModule_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	147 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_Sample/ra
      -- 
    ra_8815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3663_inst_ack_0, ack => sendModule_CP_8180_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	270 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3663_Update/ca
      -- 
    ca_8820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3663_inst_ack_1, ack => sendModule_CP_8180_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	149 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_Sample/rr
      -- 
    rr_8828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(178), ack => slice_3667_inst_req_0); -- 
    sendModule_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(149) & sendModule_CP_8180_elements(180);
      gj_sendModule_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	272 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_update_start_
      -- CP-element group 179: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_Update/cr
      -- 
    cr_8833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(179), ack => slice_3667_inst_req_1); -- 
    sendModule_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	147 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_Sample/ra
      -- 
    ra_8829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3667_inst_ack_0, ack => sendModule_CP_8180_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	270 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3667_Update/ca
      -- 
    ca_8834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3667_inst_ack_1, ack => sendModule_CP_8180_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	149 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_Sample/rr
      -- 
    rr_8842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(182), ack => slice_3671_inst_req_0); -- 
    sendModule_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(149) & sendModule_CP_8180_elements(184);
      gj_sendModule_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	272 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_update_start_
      -- CP-element group 183: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_Update/cr
      -- 
    cr_8847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(183), ack => slice_3671_inst_req_1); -- 
    sendModule_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	147 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_Sample/ra
      -- 
    ra_8843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3671_inst_ack_0, ack => sendModule_CP_8180_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	270 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3671_Update/ca
      -- 
    ca_8848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3671_inst_ack_1, ack => sendModule_CP_8180_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	149 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_Sample/rr
      -- 
    rr_8856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(186), ack => slice_3675_inst_req_0); -- 
    sendModule_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(149) & sendModule_CP_8180_elements(188);
      gj_sendModule_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	272 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_update_start_
      -- CP-element group 187: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_Update/cr
      -- 
    cr_8861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(187), ack => slice_3675_inst_req_1); -- 
    sendModule_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: 	147 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_Sample/ra
      -- 
    ra_8857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3675_inst_ack_0, ack => sendModule_CP_8180_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	270 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/slice_3675_Update/ca
      -- 
    ca_8862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3675_inst_ack_1, ack => sendModule_CP_8180_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	153 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_Sample/req
      -- 
    req_8870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(190), ack => W_output_data1_3560_delayed_14_0_3685_inst_req_0); -- 
    sendModule_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(153) & sendModule_CP_8180_elements(192);
      gj_sendModule_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	260 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_update_start_
      -- CP-element group 191: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_Update/req
      -- 
    req_8875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(191), ack => W_output_data1_3560_delayed_14_0_3685_inst_req_1); -- 
    sendModule_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: 	151 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_Sample/ack
      -- 
    ack_8871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3560_delayed_14_0_3685_inst_ack_0, ack => sendModule_CP_8180_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	258 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3687_Update/ack
      -- 
    ack_8876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3560_delayed_14_0_3685_inst_ack_1, ack => sendModule_CP_8180_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	24 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_Sample/rr
      -- 
    rr_8884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(194), ack => EQ_u2_u1_3691_inst_req_0); -- 
    sendModule_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(24) & sendModule_CP_8180_elements(196);
      gj_sendModule_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	260 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_update_start_
      -- CP-element group 195: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_Update/cr
      -- 
    cr_8889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(195), ack => EQ_u2_u1_3691_inst_req_1); -- 
    sendModule_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: 	22 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_Sample/ra
      -- 
    ra_8885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3691_inst_ack_0, ack => sendModule_CP_8180_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	258 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3691_Update/ca
      -- 
    ca_8890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3691_inst_ack_1, ack => sendModule_CP_8180_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	24 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_Sample/rr
      -- 
    rr_8898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(198), ack => EQ_u2_u1_3702_inst_req_0); -- 
    sendModule_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(24) & sendModule_CP_8180_elements(200);
      gj_sendModule_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	260 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_update_start_
      -- CP-element group 199: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_Update/cr
      -- 
    cr_8903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(199), ack => EQ_u2_u1_3702_inst_req_1); -- 
    sendModule_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: 	22 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_Sample/ra
      -- 
    ra_8899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3702_inst_ack_0, ack => sendModule_CP_8180_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	258 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3702_Update/ca
      -- 
    ca_8904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3702_inst_ack_1, ack => sendModule_CP_8180_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	153 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_Sample/req
      -- 
    req_8912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(202), ack => W_output_data1_3568_delayed_14_0_3704_inst_req_0); -- 
    sendModule_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(153) & sendModule_CP_8180_elements(204);
      gj_sendModule_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	260 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_update_start_
      -- CP-element group 203: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_Update/req
      -- 
    req_8917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(203), ack => W_output_data1_3568_delayed_14_0_3704_inst_req_1); -- 
    sendModule_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	151 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_Sample/ack
      -- 
    ack_8913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3568_delayed_14_0_3704_inst_ack_0, ack => sendModule_CP_8180_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	258 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3706_Update/ack
      -- 
    ack_8918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3568_delayed_14_0_3704_inst_ack_1, ack => sendModule_CP_8180_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	24 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_Sample/rr
      -- 
    rr_8926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(206), ack => EQ_u2_u1_3716_inst_req_0); -- 
    sendModule_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(24) & sendModule_CP_8180_elements(208);
      gj_sendModule_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	260 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_update_start_
      -- CP-element group 207: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_Update/cr
      -- 
    cr_8931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(207), ack => EQ_u2_u1_3716_inst_req_1); -- 
    sendModule_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: 	22 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_Sample/ra
      -- 
    ra_8927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3716_inst_ack_0, ack => sendModule_CP_8180_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	258 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3716_Update/ca
      -- 
    ca_8932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3716_inst_ack_1, ack => sendModule_CP_8180_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	153 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_Sample/req
      -- 
    req_8940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(210), ack => W_output_data1_3576_delayed_14_0_3718_inst_req_0); -- 
    sendModule_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(153) & sendModule_CP_8180_elements(212);
      gj_sendModule_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	260 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_update_start_
      -- CP-element group 211: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_Update/req
      -- 
    req_8945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(211), ack => W_output_data1_3576_delayed_14_0_3718_inst_req_1); -- 
    sendModule_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: 	151 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_Sample/ack
      -- 
    ack_8941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3576_delayed_14_0_3718_inst_ack_0, ack => sendModule_CP_8180_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	258 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3720_Update/ack
      -- 
    ack_8946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3576_delayed_14_0_3718_inst_ack_1, ack => sendModule_CP_8180_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	24 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_Sample/rr
      -- 
    rr_8954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(214), ack => EQ_u2_u1_3730_inst_req_0); -- 
    sendModule_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(24) & sendModule_CP_8180_elements(216);
      gj_sendModule_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	260 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_update_start_
      -- CP-element group 215: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_Update/cr
      -- 
    cr_8959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(215), ack => EQ_u2_u1_3730_inst_req_1); -- 
    sendModule_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: 	22 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_Sample/ra
      -- 
    ra_8955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3730_inst_ack_0, ack => sendModule_CP_8180_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	258 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3730_Update/ca
      -- 
    ca_8960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3730_inst_ack_1, ack => sendModule_CP_8180_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	153 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_Sample/req
      -- 
    req_8968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(218), ack => W_output_data1_3584_delayed_14_0_3732_inst_req_0); -- 
    sendModule_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(153) & sendModule_CP_8180_elements(220);
      gj_sendModule_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	260 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_update_start_
      -- CP-element group 219: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_Update/req
      -- 
    req_8973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(219), ack => W_output_data1_3584_delayed_14_0_3732_inst_req_1); -- 
    sendModule_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: 	151 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_Sample/ack
      -- 
    ack_8969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3584_delayed_14_0_3732_inst_ack_0, ack => sendModule_CP_8180_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	258 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3734_Update/ack
      -- 
    ack_8974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3584_delayed_14_0_3732_inst_ack_1, ack => sendModule_CP_8180_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	43 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_Sample/rr
      -- 
    rr_8982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(222), ack => EQ_u2_u1_3744_inst_req_0); -- 
    sendModule_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(43) & sendModule_CP_8180_elements(224);
      gj_sendModule_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	272 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_update_start_
      -- CP-element group 223: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_Update/cr
      -- 
    cr_8987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(223), ack => EQ_u2_u1_3744_inst_req_1); -- 
    sendModule_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: 	39 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_Sample/ra
      -- 
    ra_8983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3744_inst_ack_0, ack => sendModule_CP_8180_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	270 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3744_Update/ca
      -- 
    ca_8988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3744_inst_ack_1, ack => sendModule_CP_8180_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	157 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_Sample/req
      -- 
    req_8996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(226), ack => W_output_data2_3592_delayed_14_0_3746_inst_req_0); -- 
    sendModule_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(157) & sendModule_CP_8180_elements(228);
      gj_sendModule_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	272 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_update_start_
      -- CP-element group 227: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_Update/req
      -- 
    req_9001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(227), ack => W_output_data2_3592_delayed_14_0_3746_inst_req_1); -- 
    sendModule_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: 	155 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_Sample/ack
      -- 
    ack_8997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3592_delayed_14_0_3746_inst_ack_0, ack => sendModule_CP_8180_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	270 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3748_Update/ack
      -- 
    ack_9002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3592_delayed_14_0_3746_inst_ack_1, ack => sendModule_CP_8180_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	43 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_Sample/rr
      -- 
    rr_9010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(230), ack => EQ_u2_u1_3758_inst_req_0); -- 
    sendModule_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(43) & sendModule_CP_8180_elements(232);
      gj_sendModule_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	272 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	233 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_update_start_
      -- CP-element group 231: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_Update/cr
      -- 
    cr_9015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(231), ack => EQ_u2_u1_3758_inst_req_1); -- 
    sendModule_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: 	39 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_Sample/ra
      -- 
    ra_9011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3758_inst_ack_0, ack => sendModule_CP_8180_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	270 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3758_Update/ca
      -- 
    ca_9016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3758_inst_ack_1, ack => sendModule_CP_8180_elements(233)); -- 
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	157 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_Sample/req
      -- 
    req_9024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(234), ack => W_output_data2_3600_delayed_14_0_3760_inst_req_0); -- 
    sendModule_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(157) & sendModule_CP_8180_elements(236);
      gj_sendModule_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: marked-predecessors 
    -- CP-element group 235: 	272 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_update_start_
      -- CP-element group 235: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_Update/req
      -- 
    req_9029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(235), ack => W_output_data2_3600_delayed_14_0_3760_inst_req_1); -- 
    sendModule_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	155 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_Sample/ack
      -- 
    ack_9025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3600_delayed_14_0_3760_inst_ack_0, ack => sendModule_CP_8180_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	270 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3762_Update/ack
      -- 
    ack_9030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3600_delayed_14_0_3760_inst_ack_1, ack => sendModule_CP_8180_elements(237)); -- 
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	43 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_Sample/rr
      -- 
    rr_9038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(238), ack => EQ_u2_u1_3772_inst_req_0); -- 
    sendModule_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(43) & sendModule_CP_8180_elements(240);
      gj_sendModule_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: marked-predecessors 
    -- CP-element group 239: 	272 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_update_start_
      -- CP-element group 239: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_Update/cr
      -- 
    cr_9043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(239), ack => EQ_u2_u1_3772_inst_req_1); -- 
    sendModule_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: 	39 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_Sample/ra
      -- 
    ra_9039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3772_inst_ack_0, ack => sendModule_CP_8180_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	270 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3772_Update/ca
      -- 
    ca_9044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3772_inst_ack_1, ack => sendModule_CP_8180_elements(241)); -- 
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	157 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_Sample/req
      -- 
    req_9052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(242), ack => W_output_data2_3608_delayed_14_0_3774_inst_req_0); -- 
    sendModule_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(157) & sendModule_CP_8180_elements(244);
      gj_sendModule_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: marked-predecessors 
    -- CP-element group 243: 	272 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	245 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_update_start_
      -- CP-element group 243: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_Update/req
      -- 
    req_9057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(243), ack => W_output_data2_3608_delayed_14_0_3774_inst_req_1); -- 
    sendModule_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	155 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_Sample/ack
      -- 
    ack_9053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3608_delayed_14_0_3774_inst_ack_0, ack => sendModule_CP_8180_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	243 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	270 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3776_Update/ack
      -- 
    ack_9058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3608_delayed_14_0_3774_inst_ack_1, ack => sendModule_CP_8180_elements(245)); -- 
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	43 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_Sample/rr
      -- 
    rr_9066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(246), ack => EQ_u2_u1_3786_inst_req_0); -- 
    sendModule_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(43) & sendModule_CP_8180_elements(248);
      gj_sendModule_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: marked-predecessors 
    -- CP-element group 247: 	272 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_update_start_
      -- CP-element group 247: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_Update/cr
      -- 
    cr_9071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(247), ack => EQ_u2_u1_3786_inst_req_1); -- 
    sendModule_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: 	39 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_Sample/ra
      -- 
    ra_9067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3786_inst_ack_0, ack => sendModule_CP_8180_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	270 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/EQ_u2_u1_3786_Update/ca
      -- 
    ca_9072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3786_inst_ack_1, ack => sendModule_CP_8180_elements(249)); -- 
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	157 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_Sample/req
      -- 
    req_9080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(250), ack => W_output_data2_3616_delayed_14_0_3788_inst_req_0); -- 
    sendModule_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(157) & sendModule_CP_8180_elements(252);
      gj_sendModule_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: marked-predecessors 
    -- CP-element group 251: 	272 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_update_start_
      -- CP-element group 251: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_Update/req
      -- 
    req_9085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(251), ack => W_output_data2_3616_delayed_14_0_3788_inst_req_1); -- 
    sendModule_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	155 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_Sample/ack
      -- 
    ack_9081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3616_delayed_14_0_3788_inst_ack_0, ack => sendModule_CP_8180_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	270 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3790_Update/ack
      -- 
    ack_9086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3616_delayed_14_0_3788_inst_ack_1, ack => sendModule_CP_8180_elements(253)); -- 
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	134 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_Sample/req
      -- 
    req_9094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(254), ack => W_fetch_addr1_3620_delayed_8_0_3797_inst_req_0); -- 
    sendModule_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(134) & sendModule_CP_8180_elements(256);
      gj_sendModule_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: marked-predecessors 
    -- CP-element group 255: 	264 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_update_start_
      -- CP-element group 255: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_Update/req
      -- 
    req_9099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(255), ack => W_fetch_addr1_3620_delayed_8_0_3797_inst_req_1); -- 
    sendModule_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(264);
      gj_sendModule_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	129 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_Sample/ack
      -- 
    ack_9095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr1_3620_delayed_8_0_3797_inst_ack_0, ack => sendModule_CP_8180_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	262 
    -- CP-element group 257:  members (19) 
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3799_Update/ack
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_address_calculated
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_word_address_calculated
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_root_address_calculated
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_address_resized
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_addr_resize/$entry
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_addr_resize/$exit
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_addr_resize/base_resize_req
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_addr_resize/base_resize_ack
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_plus_offset/$entry
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_plus_offset/$exit
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_plus_offset/sum_rename_req
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_base_plus_offset/sum_rename_ack
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_word_addrgen/$entry
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_word_addrgen/$exit
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_word_addrgen/root_register_req
      -- CP-element group 257: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_word_addrgen/root_register_ack
      -- 
    ack_9100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr1_3620_delayed_8_0_3797_inst_ack_1, ack => sendModule_CP_8180_elements(257)); -- 
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	193 
    -- CP-element group 258: 	197 
    -- CP-element group 258: 	201 
    -- CP-element group 258: 	205 
    -- CP-element group 258: 	209 
    -- CP-element group 258: 	213 
    -- CP-element group 258: 	217 
    -- CP-element group 258: 	221 
    -- CP-element group 258: 	161 
    -- CP-element group 258: 	165 
    -- CP-element group 258: 	169 
    -- CP-element group 258: 	173 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_Sample/rr
      -- 
    rr_9108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(258), ack => CONCAT_u32_u64_3808_inst_req_0); -- 
    sendModule_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(193) & sendModule_CP_8180_elements(197) & sendModule_CP_8180_elements(201) & sendModule_CP_8180_elements(205) & sendModule_CP_8180_elements(209) & sendModule_CP_8180_elements(213) & sendModule_CP_8180_elements(217) & sendModule_CP_8180_elements(221) & sendModule_CP_8180_elements(161) & sendModule_CP_8180_elements(165) & sendModule_CP_8180_elements(169) & sendModule_CP_8180_elements(173) & sendModule_CP_8180_elements(260);
      gj_sendModule_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: marked-predecessors 
    -- CP-element group 259: 	264 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	261 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_update_start_
      -- CP-element group 259: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_Update/cr
      -- 
    cr_9113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(259), ack => CONCAT_u32_u64_3808_inst_req_1); -- 
    sendModule_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(264);
      gj_sendModule_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	191 
    -- CP-element group 260: 	195 
    -- CP-element group 260: 	199 
    -- CP-element group 260: 	203 
    -- CP-element group 260: 	207 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	211 
    -- CP-element group 260: 	215 
    -- CP-element group 260: 	219 
    -- CP-element group 260: 	159 
    -- CP-element group 260: 	163 
    -- CP-element group 260: 	167 
    -- CP-element group 260: 	171 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_Sample/ra
      -- 
    ra_9109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3808_inst_ack_0, ack => sendModule_CP_8180_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3808_Update/ca
      -- 
    ca_9114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3808_inst_ack_1, ack => sendModule_CP_8180_elements(261)); -- 
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	257 
    -- CP-element group 262: 	261 
    -- CP-element group 262: 	283 
    -- CP-element group 262: 	284 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	264 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (9) 
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/ptr_deref_3801_Split/$entry
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/ptr_deref_3801_Split/$exit
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/ptr_deref_3801_Split/split_req
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/ptr_deref_3801_Split/split_ack
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/word_access_start/$entry
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/word_access_start/word_0/$entry
      -- CP-element group 262: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/word_access_start/word_0/rr
      -- 
    rr_9152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(262), ack => ptr_deref_3801_store_0_req_0); -- 
    sendModule_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(257) & sendModule_CP_8180_elements(261) & sendModule_CP_8180_elements(283) & sendModule_CP_8180_elements(284) & sendModule_CP_8180_elements(264);
      gj_sendModule_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	265 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (5) 
      -- CP-element group 263: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_update_start_
      -- CP-element group 263: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Update/word_access_complete/$entry
      -- CP-element group 263: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Update/word_access_complete/word_0/$entry
      -- CP-element group 263: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Update/word_access_complete/word_0/cr
      -- 
    cr_9163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(263), ack => ptr_deref_3801_store_0_req_1); -- 
    sendModule_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(265);
      gj_sendModule_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	285 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	255 
    -- CP-element group 264: 	259 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (5) 
      -- CP-element group 264: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/word_access_start/$exit
      -- CP-element group 264: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/word_access_start/word_0/$exit
      -- CP-element group 264: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Sample/word_access_start/word_0/ra
      -- 
    ra_9153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3801_store_0_ack_0, ack => sendModule_CP_8180_elements(264)); -- 
    -- CP-element group 265:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	286 
    -- CP-element group 265: marked-successors 
    -- CP-element group 265: 	263 
    -- CP-element group 265:  members (5) 
      -- CP-element group 265: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Update/word_access_complete/$exit
      -- CP-element group 265: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Update/word_access_complete/word_0/$exit
      -- CP-element group 265: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_Update/word_access_complete/word_0/ca
      -- 
    ca_9164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3801_store_0_ack_1, ack => sendModule_CP_8180_elements(265)); -- 
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	141 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_Sample/req
      -- 
    req_9172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(266), ack => W_fetch_addr2_3630_delayed_8_0_3810_inst_req_0); -- 
    sendModule_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(141) & sendModule_CP_8180_elements(268);
      gj_sendModule_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	276 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_update_start_
      -- CP-element group 267: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_Update/req
      -- 
    req_9177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(267), ack => W_fetch_addr2_3630_delayed_8_0_3810_inst_req_1); -- 
    sendModule_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(276);
      gj_sendModule_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	136 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_Sample/ack
      -- 
    ack_9173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr2_3630_delayed_8_0_3810_inst_ack_0, ack => sendModule_CP_8180_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	274 
    -- CP-element group 269:  members (19) 
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/assign_stmt_3812_Update/ack
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_word_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_root_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_address_resized
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_addr_resize/$entry
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_addr_resize/$exit
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_addr_resize/base_resize_req
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_addr_resize/base_resize_ack
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_plus_offset/$entry
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_plus_offset/$exit
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_plus_offset/sum_rename_req
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_base_plus_offset/sum_rename_ack
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_word_addrgen/$entry
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_word_addrgen/$exit
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_word_addrgen/root_register_req
      -- CP-element group 269: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_word_addrgen/root_register_ack
      -- 
    ack_9178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr2_3630_delayed_8_0_3810_inst_ack_1, ack => sendModule_CP_8180_elements(269)); -- 
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	181 
    -- CP-element group 270: 	185 
    -- CP-element group 270: 	189 
    -- CP-element group 270: 	241 
    -- CP-element group 270: 	245 
    -- CP-element group 270: 	249 
    -- CP-element group 270: 	253 
    -- CP-element group 270: 	225 
    -- CP-element group 270: 	229 
    -- CP-element group 270: 	233 
    -- CP-element group 270: 	237 
    -- CP-element group 270: 	177 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_Sample/rr
      -- 
    rr_9186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(270), ack => CONCAT_u32_u64_3821_inst_req_0); -- 
    sendModule_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(181) & sendModule_CP_8180_elements(185) & sendModule_CP_8180_elements(189) & sendModule_CP_8180_elements(241) & sendModule_CP_8180_elements(245) & sendModule_CP_8180_elements(249) & sendModule_CP_8180_elements(253) & sendModule_CP_8180_elements(225) & sendModule_CP_8180_elements(229) & sendModule_CP_8180_elements(233) & sendModule_CP_8180_elements(237) & sendModule_CP_8180_elements(177) & sendModule_CP_8180_elements(272);
      gj_sendModule_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: marked-predecessors 
    -- CP-element group 271: 	276 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_update_start_
      -- CP-element group 271: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_Update/cr
      -- 
    cr_9191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(271), ack => CONCAT_u32_u64_3821_inst_req_1); -- 
    sendModule_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(276);
      gj_sendModule_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	183 
    -- CP-element group 272: 	187 
    -- CP-element group 272: 	243 
    -- CP-element group 272: 	247 
    -- CP-element group 272: 	251 
    -- CP-element group 272: 	223 
    -- CP-element group 272: 	227 
    -- CP-element group 272: 	231 
    -- CP-element group 272: 	235 
    -- CP-element group 272: 	239 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	175 
    -- CP-element group 272: 	179 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_Sample/ra
      -- 
    ra_9187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3821_inst_ack_0, ack => sendModule_CP_8180_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/CONCAT_u32_u64_3821_Update/ca
      -- 
    ca_9192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3821_inst_ack_1, ack => sendModule_CP_8180_elements(273)); -- 
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	269 
    -- CP-element group 274: 	273 
    -- CP-element group 274: 	285 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (9) 
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/ptr_deref_3814_Split/$entry
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/ptr_deref_3814_Split/$exit
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/ptr_deref_3814_Split/split_req
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/ptr_deref_3814_Split/split_ack
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/word_access_start/$entry
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/word_access_start/word_0/$entry
      -- CP-element group 274: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/word_access_start/word_0/rr
      -- 
    rr_9230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(274), ack => ptr_deref_3814_store_0_req_0); -- 
    sendModule_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(269) & sendModule_CP_8180_elements(273) & sendModule_CP_8180_elements(285) & sendModule_CP_8180_elements(276);
      gj_sendModule_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	277 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (5) 
      -- CP-element group 275: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_update_start_
      -- CP-element group 275: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Update/word_access_complete/$entry
      -- CP-element group 275: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Update/word_access_complete/word_0/$entry
      -- CP-element group 275: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Update/word_access_complete/word_0/cr
      -- 
    cr_9241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(275), ack => ptr_deref_3814_store_0_req_1); -- 
    sendModule_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(277);
      gj_sendModule_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	286 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	267 
    -- CP-element group 276: 	271 
    -- CP-element group 276: 	274 
    -- CP-element group 276: 	142 
    -- CP-element group 276: 	146 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/word_access_start/$exit
      -- CP-element group 276: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/word_access_start/word_0/$exit
      -- CP-element group 276: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Sample/word_access_start/word_0/ra
      -- CP-element group 276: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ring_reenable_memory_space_0
      -- 
    ra_9231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3814_store_0_ack_0, ack => sendModule_CP_8180_elements(276)); -- 
    -- CP-element group 277:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	286 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	275 
    -- CP-element group 277:  members (5) 
      -- CP-element group 277: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Update/word_access_complete/$exit
      -- CP-element group 277: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Update/word_access_complete/word_0/$exit
      -- CP-element group 277: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3814_Update/word_access_complete/word_0/ca
      -- 
    ca_9242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3814_store_0_ack_1, ack => sendModule_CP_8180_elements(277)); -- 
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	15 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_Sample/rr
      -- 
    rr_9250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(278), ack => SUB_u16_u16_3826_inst_req_0); -- 
    sendModule_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(15) & sendModule_CP_8180_elements(280);
      gj_sendModule_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_update_start_
      -- CP-element group 279: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_Update/cr
      -- 
    cr_9255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(279), ack => SUB_u16_u16_3826_inst_req_1); -- 
    sendModule_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_8180_elements(281);
      gj_sendModule_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	278 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_sample_completed_
      -- CP-element group 280: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_Sample/ra
      -- 
    ra_9251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3826_inst_ack_0, ack => sendModule_CP_8180_elements(280)); -- 
    -- CP-element group 281:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	16 
    -- CP-element group 281: marked-successors 
    -- CP-element group 281: 	279 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_update_completed_
      -- CP-element group 281: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/SUB_u16_u16_3826_Update/ca
      -- 
    ca_9256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3826_inst_ack_1, ack => sendModule_CP_8180_elements(281)); -- 
    -- CP-element group 282:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	15 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	16 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group sendModule_CP_8180_elements(282) is a control-delay.
    cp_element_282_delay: control_delay_element  generic map(name => " 282_delay", delay_value => 1)  port map(req => sendModule_CP_8180_elements(15), ack => sendModule_CP_8180_elements(282), clk => clk, reset =>reset);
    -- CP-element group 283:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	144 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	262 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3633_ptr_deref_3801_delay
      -- 
    -- Element group sendModule_CP_8180_elements(283) is a control-delay.
    cp_element_283_delay: control_delay_element  generic map(name => " 283_delay", delay_value => 1)  port map(req => sendModule_CP_8180_elements(144), ack => sendModule_CP_8180_elements(283), clk => clk, reset =>reset);
    -- CP-element group 284:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	148 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	262 
    -- CP-element group 284:  members (1) 
      -- CP-element group 284: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3637_ptr_deref_3801_delay
      -- 
    -- Element group sendModule_CP_8180_elements(284) is a control-delay.
    cp_element_284_delay: control_delay_element  generic map(name => " 284_delay", delay_value => 1)  port map(req => sendModule_CP_8180_elements(148), ack => sendModule_CP_8180_elements(284), clk => clk, reset =>reset);
    -- CP-element group 285:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	264 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	274 
    -- CP-element group 285:  members (1) 
      -- CP-element group 285: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/ptr_deref_3801_ptr_deref_3814_delay
      -- 
    -- Element group sendModule_CP_8180_elements(285) is a control-delay.
    cp_element_285_delay: control_delay_element  generic map(name => " 285_delay", delay_value => 1)  port map(req => sendModule_CP_8180_elements(264), ack => sendModule_CP_8180_elements(285), clk => clk, reset =>reset);
    -- CP-element group 286:  join  transition  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	18 
    -- CP-element group 286: 	123 
    -- CP-element group 286: 	127 
    -- CP-element group 286: 	131 
    -- CP-element group 286: 	265 
    -- CP-element group 286: 	276 
    -- CP-element group 286: 	277 
    -- CP-element group 286: 	138 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	12 
    -- CP-element group 286:  members (1) 
      -- CP-element group 286: 	 branch_block_stmt_3479/do_while_stmt_3495/do_while_stmt_3495_loop_body/$exit
      -- 
    sendModule_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_8180_elements(18) & sendModule_CP_8180_elements(123) & sendModule_CP_8180_elements(127) & sendModule_CP_8180_elements(131) & sendModule_CP_8180_elements(265) & sendModule_CP_8180_elements(276) & sendModule_CP_8180_elements(277) & sendModule_CP_8180_elements(138);
      gj_sendModule_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_8180_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	11 
    -- CP-element group 287: successors 
    -- CP-element group 287:  members (2) 
      -- CP-element group 287: 	 branch_block_stmt_3479/do_while_stmt_3495/loop_exit/$exit
      -- CP-element group 287: 	 branch_block_stmt_3479/do_while_stmt_3495/loop_exit/ack
      -- 
    ack_9265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3495_branch_ack_0, ack => sendModule_CP_8180_elements(287)); -- 
    -- CP-element group 288:  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	11 
    -- CP-element group 288: successors 
    -- CP-element group 288:  members (2) 
      -- CP-element group 288: 	 branch_block_stmt_3479/do_while_stmt_3495/loop_taken/$exit
      -- CP-element group 288: 	 branch_block_stmt_3479/do_while_stmt_3495/loop_taken/ack
      -- 
    ack_9269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3495_branch_ack_1, ack => sendModule_CP_8180_elements(288)); -- 
    -- CP-element group 289:  transition  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	9 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	1 
    -- CP-element group 289:  members (1) 
      -- CP-element group 289: 	 branch_block_stmt_3479/do_while_stmt_3495/$exit
      -- 
    sendModule_CP_8180_elements(289) <= sendModule_CP_8180_elements(9);
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	1 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_update_start_
      -- CP-element group 290: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_Sample/ack
      -- CP-element group 290: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_Update/req
      -- 
    ack_9282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3838_inst_ack_0, ack => sendModule_CP_8180_elements(290)); -- 
    req_9286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_8180_elements(290), ack => WPIPE_input_done_pipe_3838_inst_req_1); -- 
    -- CP-element group 291:  transition  place  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (8) 
      -- CP-element group 291: 	 $exit
      -- CP-element group 291: 	 branch_block_stmt_3479/$exit
      -- CP-element group 291: 	 branch_block_stmt_3479/branch_block_stmt_3479__exit__
      -- CP-element group 291: 	 branch_block_stmt_3479/assign_stmt_3840__exit__
      -- CP-element group 291: 	 branch_block_stmt_3479/assign_stmt_3840/$exit
      -- CP-element group 291: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_Update/$exit
      -- CP-element group 291: 	 branch_block_stmt_3479/assign_stmt_3840/WPIPE_input_done_pipe_3838_Update/ack
      -- 
    ack_9287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3838_inst_ack_1, ack => sendModule_CP_8180_elements(291)); -- 
    sendModule_do_while_stmt_3495_terminator_9270: loop_terminator -- 
      generic map (name => " sendModule_do_while_stmt_3495_terminator_9270", max_iterations_in_flight =>15) 
      port map(loop_body_exit => sendModule_CP_8180_elements(12),loop_continue => sendModule_CP_8180_elements(288),loop_terminate => sendModule_CP_8180_elements(287),loop_back => sendModule_CP_8180_elements(10),loop_exit => sendModule_CP_8180_elements(9),clk => clk, reset => reset); -- 
    phi_stmt_3497_phi_seq_8302_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_8180_elements(27);
      sendModule_CP_8180_elements(30)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_8180_elements(30);
      sendModule_CP_8180_elements(31)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_8180_elements(32);
      sendModule_CP_8180_elements(28) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_8180_elements(25);
      sendModule_CP_8180_elements(34)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_8180_elements(36);
      sendModule_CP_8180_elements(35)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_8180_elements(37);
      sendModule_CP_8180_elements(26) <= phi_mux_reqs(1);
      phi_stmt_3497_phi_seq_8302 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3497_phi_seq_8302") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_8180_elements(17), 
          phi_sample_ack => sendModule_CP_8180_elements(23), 
          phi_update_req => sendModule_CP_8180_elements(19), 
          phi_update_ack => sendModule_CP_8180_elements(24), 
          phi_mux_ack => sendModule_CP_8180_elements(29), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3502_phi_seq_8356_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_8180_elements(46);
      sendModule_CP_8180_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_8180_elements(53);
      sendModule_CP_8180_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_8180_elements(54);
      sendModule_CP_8180_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_8180_elements(44);
      sendModule_CP_8180_elements(55)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_8180_elements(57);
      sendModule_CP_8180_elements(56)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_8180_elements(58);
      sendModule_CP_8180_elements(45) <= phi_mux_reqs(1);
      phi_stmt_3502_phi_seq_8356 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3502_phi_seq_8356") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_8180_elements(40), 
          phi_sample_ack => sendModule_CP_8180_elements(41), 
          phi_update_req => sendModule_CP_8180_elements(42), 
          phi_update_ack => sendModule_CP_8180_elements(43), 
          phi_mux_ack => sendModule_CP_8180_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3507_phi_seq_8400_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_8180_elements(67);
      sendModule_CP_8180_elements(70)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_8180_elements(70);
      sendModule_CP_8180_elements(71)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_8180_elements(72);
      sendModule_CP_8180_elements(68) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_8180_elements(65);
      sendModule_CP_8180_elements(74)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_8180_elements(76);
      sendModule_CP_8180_elements(75)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_8180_elements(77);
      sendModule_CP_8180_elements(66) <= phi_mux_reqs(1);
      phi_stmt_3507_phi_seq_8400 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3507_phi_seq_8400") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_8180_elements(61), 
          phi_sample_ack => sendModule_CP_8180_elements(62), 
          phi_update_req => sendModule_CP_8180_elements(63), 
          phi_update_ack => sendModule_CP_8180_elements(64), 
          phi_mux_ack => sendModule_CP_8180_elements(69), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3512_phi_seq_8444_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_8180_elements(86);
      sendModule_CP_8180_elements(89)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_8180_elements(89);
      sendModule_CP_8180_elements(90)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_8180_elements(91);
      sendModule_CP_8180_elements(87) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_8180_elements(84);
      sendModule_CP_8180_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_8180_elements(95);
      sendModule_CP_8180_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_8180_elements(96);
      sendModule_CP_8180_elements(85) <= phi_mux_reqs(1);
      phi_stmt_3512_phi_seq_8444 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3512_phi_seq_8444") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_8180_elements(80), 
          phi_sample_ack => sendModule_CP_8180_elements(81), 
          phi_update_req => sendModule_CP_8180_elements(82), 
          phi_update_ack => sendModule_CP_8180_elements(83), 
          phi_mux_ack => sendModule_CP_8180_elements(88), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3517_phi_seq_8488_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_8180_elements(105);
      sendModule_CP_8180_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_8180_elements(108);
      sendModule_CP_8180_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_8180_elements(110);
      sendModule_CP_8180_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_8180_elements(103);
      sendModule_CP_8180_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_8180_elements(114);
      sendModule_CP_8180_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_8180_elements(115);
      sendModule_CP_8180_elements(104) <= phi_mux_reqs(1);
      phi_stmt_3517_phi_seq_8488 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3517_phi_seq_8488") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_8180_elements(99), 
          phi_sample_ack => sendModule_CP_8180_elements(100), 
          phi_update_req => sendModule_CP_8180_elements(101), 
          phi_update_ack => sendModule_CP_8180_elements(102), 
          phi_mux_ack => sendModule_CP_8180_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_8254_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= sendModule_CP_8180_elements(13);
        preds(1)  <= sendModule_CP_8180_elements(14);
        entry_tmerge_8254 : transition_merge -- 
          generic map(name => " entry_tmerge_8254")
          port map (preds => preds, symbol_out => sendModule_CP_8180_elements(15));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_3545_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3554_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3563_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_3592_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3602_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3606_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3804_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3807_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3817_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3820_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_3808_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_3821_wire : std_logic_vector(63 downto 0);
    signal EQ_u2_u1_3559_3559_delayed_14_0_3692 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3567_3567_delayed_14_0_3703 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3575_3575_delayed_14_0_3717 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3583_3583_delayed_14_0_3731 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3591_3591_delayed_14_0_3745 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3599_3599_delayed_14_0_3759 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3607_3607_delayed_14_0_3773 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3615_3615_delayed_14_0_3787 : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_3616_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_3626_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_3492_wire : std_logic_vector(15 downto 0);
    signal MUX_3556_wire : std_logic_vector(15 downto 0);
    signal MUX_3594_wire : std_logic_vector(31 downto 0);
    signal MUX_3608_wire : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_3833_wire : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_3413_3413_delayed_1_0_3532 : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_3644_3644_delayed_1_0_3827 : std_logic_vector(15 downto 0);
    signal UGE_u16_u1_3537_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_3831_wire : std_logic_vector(0 downto 0);
    signal address1_3497 : std_logic_vector(31 downto 0);
    signal address2_3502 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3618_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3618_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3618_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3618_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3618_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3618_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3628_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3628_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3628_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3628_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3628_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3628_root_address : std_logic_vector(13 downto 0);
    signal cb_3485 : std_logic_vector(15 downto 0);
    signal chl_3507 : std_logic_vector(15 downto 0);
    signal chl_change_3539 : std_logic_vector(0 downto 0);
    signal chl_out_3488 : std_logic_vector(15 downto 0);
    signal col_3512 : std_logic_vector(15 downto 0);
    signal continue_flag_3835 : std_logic_vector(0 downto 0);
    signal fetch_addr1_3620 : std_logic_vector(31 downto 0);
    signal fetch_addr1_3620_delayed_8_0_3799 : std_logic_vector(31 downto 0);
    signal fetch_addr2_3630 : std_logic_vector(31 downto 0);
    signal fetch_addr2_3630_delayed_8_0_3812 : std_logic_vector(31 downto 0);
    signal fetch_val1_3634 : std_logic_vector(63 downto 0);
    signal fetch_val2_3638 : std_logic_vector(63 downto 0);
    signal konst_3530_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3542_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3544_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3550_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3553_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3562_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3615_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3625_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3690_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3701_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3715_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3729_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3743_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3757_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3771_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3785_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3825_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3839_wire_constant : std_logic_vector(7 downto 0);
    signal location1_3680 : std_logic_vector(1 downto 0);
    signal location2_3684 : std_logic_vector(1 downto 0);
    signal n_address1_3596 : std_logic_vector(31 downto 0);
    signal n_address1_3596_3501_buffered : std_logic_vector(31 downto 0);
    signal n_address2_3610 : std_logic_vector(31 downto 0);
    signal n_address2_3610_3506_buffered : std_logic_vector(31 downto 0);
    signal n_chl_3566 : std_logic_vector(15 downto 0);
    signal n_chl_3566_3511_buffered : std_logic_vector(15 downto 0);
    signal n_col_3547 : std_logic_vector(15 downto 0);
    signal n_col_3547_3516_buffered : std_logic_vector(15 downto 0);
    signal n_row_3558 : std_logic_vector(15 downto 0);
    signal n_row_3558_3521_buffered : std_logic_vector(15 downto 0);
    signal output_data1_3560_delayed_14_0_3687 : std_logic_vector(15 downto 0);
    signal output_data1_3568_delayed_14_0_3706 : std_logic_vector(15 downto 0);
    signal output_data1_3576_delayed_14_0_3720 : std_logic_vector(15 downto 0);
    signal output_data1_3584_delayed_14_0_3734 : std_logic_vector(15 downto 0);
    signal output_data1_3641 : std_logic_vector(15 downto 0);
    signal output_data2_3592_delayed_14_0_3748 : std_logic_vector(15 downto 0);
    signal output_data2_3600_delayed_14_0_3762 : std_logic_vector(15 downto 0);
    signal output_data2_3608_delayed_14_0_3776 : std_logic_vector(15 downto 0);
    signal output_data2_3616_delayed_14_0_3790 : std_logic_vector(15 downto 0);
    signal output_data2_3644 : std_logic_vector(15 downto 0);
    signal ptr_deref_3633_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3633_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3633_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3633_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3633_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3637_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3637_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3637_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3637_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3637_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3801_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3801_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3801_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3801_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3801_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3801_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3814_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3814_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3814_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3814_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3814_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3814_word_offset_0 : std_logic_vector(13 downto 0);
    signal rb_3482 : std_logic_vector(15 downto 0);
    signal row_3517 : std_logic_vector(15 downto 0);
    signal row_change_3527 : std_logic_vector(0 downto 0);
    signal row_size_3494 : std_logic_vector(31 downto 0);
    signal tmp1_3575 : std_logic_vector(31 downto 0);
    signal tmp2_3584 : std_logic_vector(31 downto 0);
    signal type_cast_3447_3447_delayed_1_0_3570 : std_logic_vector(31 downto 0);
    signal type_cast_3453_3453_delayed_1_0_3579 : std_logic_vector(31 downto 0);
    signal type_cast_3500_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3505_wire : std_logic_vector(31 downto 0);
    signal type_cast_3510_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3515_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3520_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3588_wire : std_logic_vector(31 downto 0);
    signal type_cast_3600_wire : std_logic_vector(31 downto 0);
    signal type_cast_3617_resized : std_logic_vector(13 downto 0);
    signal type_cast_3617_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3617_wire : std_logic_vector(63 downto 0);
    signal type_cast_3627_resized : std_logic_vector(13 downto 0);
    signal type_cast_3627_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3627_wire : std_logic_vector(63 downto 0);
    signal w11_3648 : std_logic_vector(15 downto 0);
    signal w12_3652 : std_logic_vector(15 downto 0);
    signal w13_3656 : std_logic_vector(15 downto 0);
    signal w14_3660 : std_logic_vector(15 downto 0);
    signal w21_3664 : std_logic_vector(15 downto 0);
    signal w22_3668 : std_logic_vector(15 downto 0);
    signal w23_3672 : std_logic_vector(15 downto 0);
    signal w24_3676 : std_logic_vector(15 downto 0);
    signal wb11_3698 : std_logic_vector(15 downto 0);
    signal wb12_3712 : std_logic_vector(15 downto 0);
    signal wb13_3726 : std_logic_vector(15 downto 0);
    signal wb14_3740 : std_logic_vector(15 downto 0);
    signal wb21_3754 : std_logic_vector(15 downto 0);
    signal wb22_3768 : std_logic_vector(15 downto 0);
    signal wb23_3782 : std_logic_vector(15 downto 0);
    signal wb24_3796 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_3618_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3618_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3618_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3618_resized_base_address <= "00000000000000";
    array_obj_ref_3628_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3628_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3628_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3628_resized_base_address <= "00000000000000";
    konst_3530_wire_constant <= "0000000000000001";
    konst_3542_wire_constant <= "0000000000000001";
    konst_3544_wire_constant <= "0000000000000001";
    konst_3550_wire_constant <= "0000000000000001";
    konst_3553_wire_constant <= "0000000000000010";
    konst_3562_wire_constant <= "0000000000000001";
    konst_3615_wire_constant <= "00000000000000000000000000000010";
    konst_3625_wire_constant <= "00000000000000000000000000000010";
    konst_3690_wire_constant <= "00";
    konst_3701_wire_constant <= "01";
    konst_3715_wire_constant <= "10";
    konst_3729_wire_constant <= "11";
    konst_3743_wire_constant <= "00";
    konst_3757_wire_constant <= "01";
    konst_3771_wire_constant <= "10";
    konst_3785_wire_constant <= "11";
    konst_3825_wire_constant <= "0000000000000001";
    konst_3839_wire_constant <= "00000001";
    ptr_deref_3633_word_offset_0 <= "00000000000000";
    ptr_deref_3637_word_offset_0 <= "00000000000000";
    ptr_deref_3801_word_offset_0 <= "00000000000000";
    ptr_deref_3814_word_offset_0 <= "00000000000000";
    type_cast_3500_wire_constant <= "00000000000000000000000000000000";
    type_cast_3510_wire_constant <= "0000000000000000";
    type_cast_3515_wire_constant <= "0000000000000001";
    type_cast_3520_wire_constant <= "0000000000000001";
    phi_stmt_3497: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3500_wire_constant & n_address1_3596_3501_buffered;
      req <= phi_stmt_3497_req_0 & phi_stmt_3497_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3497",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3497_ack_0,
          idata => idata,
          odata => address1_3497,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3497
    phi_stmt_3502: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3505_wire & n_address2_3610_3506_buffered;
      req <= phi_stmt_3502_req_0 & phi_stmt_3502_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3502",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3502_ack_0,
          idata => idata,
          odata => address2_3502,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3502
    phi_stmt_3507: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3510_wire_constant & n_chl_3566_3511_buffered;
      req <= phi_stmt_3507_req_0 & phi_stmt_3507_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3507",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3507_ack_0,
          idata => idata,
          odata => chl_3507,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3507
    phi_stmt_3512: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3515_wire_constant & n_col_3547_3516_buffered;
      req <= phi_stmt_3512_req_0 & phi_stmt_3512_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3512",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3512_ack_0,
          idata => idata,
          odata => col_3512,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3512
    phi_stmt_3517: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3520_wire_constant & n_row_3558_3521_buffered;
      req <= phi_stmt_3517_req_0 & phi_stmt_3517_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3517",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3517_ack_0,
          idata => idata,
          odata => row_3517,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3517
    -- flow-through select operator MUX_3546_inst
    n_col_3547 <= konst_3542_wire_constant when (row_change_3527(0) /=  '0') else ADD_u16_u16_3545_wire;
    -- flow-through select operator MUX_3556_inst
    MUX_3556_wire <= ADD_u16_u16_3554_wire when (row_change_3527(0) /=  '0') else row_3517;
    -- flow-through select operator MUX_3557_inst
    n_row_3558 <= konst_3550_wire_constant when (chl_change_3539(0) /=  '0') else MUX_3556_wire;
    -- flow-through select operator MUX_3565_inst
    n_chl_3566 <= ADD_u16_u16_3563_wire when (chl_change_3539(0) /=  '0') else chl_3507;
    -- flow-through select operator MUX_3594_inst
    MUX_3594_wire <= ADD_u32_u32_3592_wire when (row_change_3527(0) /=  '0') else tmp1_3575;
    -- flow-through select operator MUX_3595_inst
    n_address1_3596 <= type_cast_3588_wire when (chl_change_3539(0) /=  '0') else MUX_3594_wire;
    -- flow-through select operator MUX_3608_inst
    MUX_3608_wire <= ADD_u32_u32_3606_wire when (row_change_3527(0) /=  '0') else tmp2_3584;
    -- flow-through select operator MUX_3609_inst
    n_address2_3610 <= ADD_u32_u32_3602_wire when (chl_change_3539(0) /=  '0') else MUX_3608_wire;
    -- flow-through select operator MUX_3697_inst
    wb11_3698 <= output_data1_3560_delayed_14_0_3687 when (EQ_u2_u1_3559_3559_delayed_14_0_3692(0) /=  '0') else w11_3648;
    -- flow-through select operator MUX_3711_inst
    wb12_3712 <= output_data1_3568_delayed_14_0_3706 when (EQ_u2_u1_3567_3567_delayed_14_0_3703(0) /=  '0') else w12_3652;
    -- flow-through select operator MUX_3725_inst
    wb13_3726 <= output_data1_3576_delayed_14_0_3720 when (EQ_u2_u1_3575_3575_delayed_14_0_3717(0) /=  '0') else w13_3656;
    -- flow-through select operator MUX_3739_inst
    wb14_3740 <= output_data1_3584_delayed_14_0_3734 when (EQ_u2_u1_3583_3583_delayed_14_0_3731(0) /=  '0') else w14_3660;
    -- flow-through select operator MUX_3753_inst
    wb21_3754 <= output_data2_3592_delayed_14_0_3748 when (EQ_u2_u1_3591_3591_delayed_14_0_3745(0) /=  '0') else w21_3664;
    -- flow-through select operator MUX_3767_inst
    wb22_3768 <= output_data2_3600_delayed_14_0_3762 when (EQ_u2_u1_3599_3599_delayed_14_0_3759(0) /=  '0') else w22_3668;
    -- flow-through select operator MUX_3781_inst
    wb23_3782 <= output_data2_3608_delayed_14_0_3776 when (EQ_u2_u1_3607_3607_delayed_14_0_3773(0) /=  '0') else w23_3672;
    -- flow-through select operator MUX_3795_inst
    wb24_3796 <= output_data2_3616_delayed_14_0_3790 when (EQ_u2_u1_3615_3615_delayed_14_0_3787(0) /=  '0') else w24_3676;
    slice_3647_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3647_inst_req_0;
      slice_3647_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3647_inst_req_1;
      slice_3647_inst_ack_1<= update_ack(0);
      slice_3647_inst: SliceSplitProtocol generic map(name => "slice_3647_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3634, dout => w11_3648, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3651_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3651_inst_req_0;
      slice_3651_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3651_inst_req_1;
      slice_3651_inst_ack_1<= update_ack(0);
      slice_3651_inst: SliceSplitProtocol generic map(name => "slice_3651_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3634, dout => w12_3652, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3655_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3655_inst_req_0;
      slice_3655_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3655_inst_req_1;
      slice_3655_inst_ack_1<= update_ack(0);
      slice_3655_inst: SliceSplitProtocol generic map(name => "slice_3655_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3634, dout => w13_3656, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3659_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3659_inst_req_0;
      slice_3659_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3659_inst_req_1;
      slice_3659_inst_ack_1<= update_ack(0);
      slice_3659_inst: SliceSplitProtocol generic map(name => "slice_3659_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3634, dout => w14_3660, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3663_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3663_inst_req_0;
      slice_3663_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3663_inst_req_1;
      slice_3663_inst_ack_1<= update_ack(0);
      slice_3663_inst: SliceSplitProtocol generic map(name => "slice_3663_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3638, dout => w21_3664, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3667_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3667_inst_req_0;
      slice_3667_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3667_inst_req_1;
      slice_3667_inst_ack_1<= update_ack(0);
      slice_3667_inst: SliceSplitProtocol generic map(name => "slice_3667_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3638, dout => w22_3668, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3671_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3671_inst_req_0;
      slice_3671_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3671_inst_req_1;
      slice_3671_inst_ack_1<= update_ack(0);
      slice_3671_inst: SliceSplitProtocol generic map(name => "slice_3671_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3638, dout => w23_3672, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3675_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3675_inst_req_0;
      slice_3675_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3675_inst_req_1;
      slice_3675_inst_ack_1<= update_ack(0);
      slice_3675_inst: SliceSplitProtocol generic map(name => "slice_3675_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3638, dout => w24_3676, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_fetch_addr1_3620_delayed_8_0_3797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr1_3620_delayed_8_0_3797_inst_req_0;
      W_fetch_addr1_3620_delayed_8_0_3797_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr1_3620_delayed_8_0_3797_inst_req_1;
      W_fetch_addr1_3620_delayed_8_0_3797_inst_ack_1<= rack(0);
      W_fetch_addr1_3620_delayed_8_0_3797_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr1_3620_delayed_8_0_3797_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr1_3620,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_3620_delayed_8_0_3799,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_addr2_3630_delayed_8_0_3810_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr2_3630_delayed_8_0_3810_inst_req_0;
      W_fetch_addr2_3630_delayed_8_0_3810_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr2_3630_delayed_8_0_3810_inst_req_1;
      W_fetch_addr2_3630_delayed_8_0_3810_inst_ack_1<= rack(0);
      W_fetch_addr2_3630_delayed_8_0_3810_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr2_3630_delayed_8_0_3810_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr2_3630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_3630_delayed_8_0_3812,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3560_delayed_14_0_3685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3560_delayed_14_0_3685_inst_req_0;
      W_output_data1_3560_delayed_14_0_3685_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3560_delayed_14_0_3685_inst_req_1;
      W_output_data1_3560_delayed_14_0_3685_inst_ack_1<= rack(0);
      W_output_data1_3560_delayed_14_0_3685_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3560_delayed_14_0_3685_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3560_delayed_14_0_3687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3568_delayed_14_0_3704_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3568_delayed_14_0_3704_inst_req_0;
      W_output_data1_3568_delayed_14_0_3704_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3568_delayed_14_0_3704_inst_req_1;
      W_output_data1_3568_delayed_14_0_3704_inst_ack_1<= rack(0);
      W_output_data1_3568_delayed_14_0_3704_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3568_delayed_14_0_3704_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3568_delayed_14_0_3706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3576_delayed_14_0_3718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3576_delayed_14_0_3718_inst_req_0;
      W_output_data1_3576_delayed_14_0_3718_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3576_delayed_14_0_3718_inst_req_1;
      W_output_data1_3576_delayed_14_0_3718_inst_ack_1<= rack(0);
      W_output_data1_3576_delayed_14_0_3718_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3576_delayed_14_0_3718_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3576_delayed_14_0_3720,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3584_delayed_14_0_3732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3584_delayed_14_0_3732_inst_req_0;
      W_output_data1_3584_delayed_14_0_3732_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3584_delayed_14_0_3732_inst_req_1;
      W_output_data1_3584_delayed_14_0_3732_inst_ack_1<= rack(0);
      W_output_data1_3584_delayed_14_0_3732_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3584_delayed_14_0_3732_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3584_delayed_14_0_3734,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3592_delayed_14_0_3746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3592_delayed_14_0_3746_inst_req_0;
      W_output_data2_3592_delayed_14_0_3746_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3592_delayed_14_0_3746_inst_req_1;
      W_output_data2_3592_delayed_14_0_3746_inst_ack_1<= rack(0);
      W_output_data2_3592_delayed_14_0_3746_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3592_delayed_14_0_3746_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3592_delayed_14_0_3748,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3600_delayed_14_0_3760_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3600_delayed_14_0_3760_inst_req_0;
      W_output_data2_3600_delayed_14_0_3760_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3600_delayed_14_0_3760_inst_req_1;
      W_output_data2_3600_delayed_14_0_3760_inst_ack_1<= rack(0);
      W_output_data2_3600_delayed_14_0_3760_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3600_delayed_14_0_3760_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3600_delayed_14_0_3762,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3608_delayed_14_0_3774_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3608_delayed_14_0_3774_inst_req_0;
      W_output_data2_3608_delayed_14_0_3774_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3608_delayed_14_0_3774_inst_req_1;
      W_output_data2_3608_delayed_14_0_3774_inst_ack_1<= rack(0);
      W_output_data2_3608_delayed_14_0_3774_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3608_delayed_14_0_3774_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3608_delayed_14_0_3776,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3616_delayed_14_0_3788_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3616_delayed_14_0_3788_inst_req_0;
      W_output_data2_3616_delayed_14_0_3788_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3616_delayed_14_0_3788_inst_req_1;
      W_output_data2_3616_delayed_14_0_3788_inst_ack_1<= rack(0);
      W_output_data2_3616_delayed_14_0_3788_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3616_delayed_14_0_3788_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3616_delayed_14_0_3790,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3619_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3619_final_reg_req_0;
      addr_of_3619_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3619_final_reg_req_1;
      addr_of_3619_final_reg_ack_1<= rack(0);
      addr_of_3619_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3619_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3618_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_3620,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3629_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3629_final_reg_req_0;
      addr_of_3629_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3629_final_reg_req_1;
      addr_of_3629_final_reg_ack_1<= rack(0);
      addr_of_3629_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3629_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3628_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_3630,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_3596_3501_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_3596_3501_buf_req_0;
      n_address1_3596_3501_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_3596_3501_buf_req_1;
      n_address1_3596_3501_buf_ack_1<= rack(0);
      n_address1_3596_3501_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_3596_3501_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_3596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_3596_3501_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_3610_3506_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_3610_3506_buf_req_0;
      n_address2_3610_3506_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_3610_3506_buf_req_1;
      n_address2_3610_3506_buf_ack_1<= rack(0);
      n_address2_3610_3506_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_3610_3506_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_3610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_3610_3506_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_3566_3511_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_3566_3511_buf_req_0;
      n_chl_3566_3511_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_3566_3511_buf_req_1;
      n_chl_3566_3511_buf_ack_1<= rack(0);
      n_chl_3566_3511_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_3566_3511_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_3566,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_3566_3511_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_3547_3516_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_3547_3516_buf_req_0;
      n_col_3547_3516_buf_ack_0<= wack(0);
      rreq(0) <= n_col_3547_3516_buf_req_1;
      n_col_3547_3516_buf_ack_1<= rack(0);
      n_col_3547_3516_buf : InterlockBuffer generic map ( -- 
        name => "n_col_3547_3516_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_3547,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_3547_3516_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_3558_3521_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_3558_3521_buf_req_0;
      n_row_3558_3521_buf_ack_0<= wack(0);
      rreq(0) <= n_row_3558_3521_buf_req_1;
      n_row_3558_3521_buf_ack_1<= rack(0);
      n_row_3558_3521_buf : InterlockBuffer generic map ( -- 
        name => "n_row_3558_3521_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_3558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_3558_3521_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3493_inst
    process(MUL_u16_u16_3492_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_3492_wire(15 downto 0);
      row_size_3494 <= tmp_var; -- 
    end process;
    type_cast_3505_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3505_inst_req_0;
      type_cast_3505_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3505_inst_req_1;
      type_cast_3505_inst_ack_1<= rack(0);
      type_cast_3505_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3505_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => row_size_3494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3505_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3569_inst_req_0;
      type_cast_3569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3569_inst_req_1;
      type_cast_3569_inst_ack_1<= rack(0);
      type_cast_3569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3569_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_3488,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3447_3447_delayed_1_0_3570,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3578_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3578_inst_req_0;
      type_cast_3578_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3578_inst_req_1;
      type_cast_3578_inst_ack_1<= rack(0);
      type_cast_3578_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3578_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_3488,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3453_3453_delayed_1_0_3579,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3588_inst
    process(n_chl_3566) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3566(15 downto 0);
      type_cast_3588_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3600_inst
    process(n_chl_3566) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3566(15 downto 0);
      type_cast_3600_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3617_inst
    process(LSHR_u32_u32_3616_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3616_wire(31 downto 0);
      type_cast_3617_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3627_inst
    process(LSHR_u32_u32_3626_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3626_wire(31 downto 0);
      type_cast_3627_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3679_inst
    process(address1_3497) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := address1_3497(1 downto 0);
      location1_3680 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3683_inst
    process(address2_3502) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := address2_3502(1 downto 0);
      location2_3684 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_3618_index_1_rename
    process(type_cast_3617_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3617_resized;
      ov(13 downto 0) := iv;
      type_cast_3617_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3618_index_1_resize
    process(type_cast_3617_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3617_wire;
      ov := iv(13 downto 0);
      type_cast_3617_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3618_root_address_inst
    process(array_obj_ref_3618_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3618_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3618_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3628_index_1_rename
    process(type_cast_3627_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3627_resized;
      ov(13 downto 0) := iv;
      type_cast_3627_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3628_index_1_resize
    process(type_cast_3627_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3627_wire;
      ov := iv(13 downto 0);
      type_cast_3627_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3628_root_address_inst
    process(array_obj_ref_3628_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3628_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3628_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3633_addr_0
    process(ptr_deref_3633_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3633_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3633_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3633_base_resize
    process(fetch_addr1_3620) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_3620;
      ov := iv(13 downto 0);
      ptr_deref_3633_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3633_gather_scatter
    process(ptr_deref_3633_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3633_data_0;
      ov(63 downto 0) := iv;
      fetch_val1_3634 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3633_root_address_inst
    process(ptr_deref_3633_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3633_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3633_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3637_addr_0
    process(ptr_deref_3637_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3637_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3637_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3637_base_resize
    process(fetch_addr2_3630) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_3630;
      ov := iv(13 downto 0);
      ptr_deref_3637_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3637_gather_scatter
    process(ptr_deref_3637_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3637_data_0;
      ov(63 downto 0) := iv;
      fetch_val2_3638 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3637_root_address_inst
    process(ptr_deref_3637_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3637_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3637_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3801_addr_0
    process(ptr_deref_3801_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3801_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3801_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3801_base_resize
    process(fetch_addr1_3620_delayed_8_0_3799) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_3620_delayed_8_0_3799;
      ov := iv(13 downto 0);
      ptr_deref_3801_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3801_gather_scatter
    process(CONCAT_u32_u64_3808_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3808_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3801_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3801_root_address_inst
    process(ptr_deref_3801_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3801_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3801_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3814_addr_0
    process(ptr_deref_3814_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3814_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3814_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3814_base_resize
    process(fetch_addr2_3630_delayed_8_0_3812) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_3630_delayed_8_0_3812;
      ov := iv(13 downto 0);
      ptr_deref_3814_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3814_gather_scatter
    process(CONCAT_u32_u64_3821_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3821_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3814_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3814_root_address_inst
    process(ptr_deref_3814_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3814_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3814_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_3495_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_3835;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3495_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3495_branch_req_0,
          ack0 => do_while_stmt_3495_branch_ack_0,
          ack1 => do_while_stmt_3495_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3545_inst
    process(col_3512) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_3512, konst_3544_wire_constant, tmp_var);
      ADD_u16_u16_3545_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3554_inst
    process(row_3517) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_3517, konst_3553_wire_constant, tmp_var);
      ADD_u16_u16_3554_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3563_inst
    process(chl_3507) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_3507, konst_3562_wire_constant, tmp_var);
      ADD_u16_u16_3563_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3574_inst
    process(address1_3497, type_cast_3447_3447_delayed_1_0_3570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_3497, type_cast_3447_3447_delayed_1_0_3570, tmp_var);
      tmp1_3575 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3583_inst
    process(address2_3502, type_cast_3453_3453_delayed_1_0_3579) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_3502, type_cast_3453_3453_delayed_1_0_3579, tmp_var);
      tmp2_3584 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3592_inst
    process(tmp1_3575, row_size_3494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_3575, row_size_3494, tmp_var);
      ADD_u32_u32_3592_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3602_inst
    process(type_cast_3600_wire, row_size_3494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_3600_wire, row_size_3494, tmp_var);
      ADD_u32_u32_3602_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3606_inst
    process(tmp2_3584, row_size_3494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_3584, row_size_3494, tmp_var);
      ADD_u32_u32_3606_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3538_inst
    process(row_change_3527, UGE_u16_u1_3537_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(row_change_3527, UGE_u16_u1_3537_wire, tmp_var);
      chl_change_3539 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3804_inst
    process(wb11_3698, wb12_3712) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb11_3698, wb12_3712, tmp_var);
      CONCAT_u16_u32_3804_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3807_inst
    process(wb13_3726, wb14_3740) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb13_3726, wb14_3740, tmp_var);
      CONCAT_u16_u32_3807_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3817_inst
    process(wb21_3754, wb22_3768) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb21_3754, wb22_3768, tmp_var);
      CONCAT_u16_u32_3817_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3820_inst
    process(wb23_3782, wb24_3796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb23_3782, wb24_3796, tmp_var);
      CONCAT_u16_u32_3820_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : CONCAT_u32_u64_3808_inst 
    ApConcat_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3804_wire & CONCAT_u16_u32_3807_wire;
      CONCAT_u32_u64_3808_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3808_inst_req_0;
      CONCAT_u32_u64_3808_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3808_inst_req_1;
      CONCAT_u32_u64_3808_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_13_gI: SplitGuardInterface generic map(name => "ApConcat_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : CONCAT_u32_u64_3821_inst 
    ApConcat_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3817_wire & CONCAT_u16_u32_3820_wire;
      CONCAT_u32_u64_3821_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3821_inst_req_0;
      CONCAT_u32_u64_3821_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3821_inst_req_1;
      CONCAT_u32_u64_3821_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_14_gI: SplitGuardInterface generic map(name => "ApConcat_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- binary operator EQ_u16_u1_3526_inst
    process(col_3512, cb_3485) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_3512, cb_3485, tmp_var);
      row_change_3527 <= tmp_var; --
    end process;
    -- shared split operator group (16) : EQ_u2_u1_3691_inst 
    ApIntEq_group_16: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3680;
      EQ_u2_u1_3559_3559_delayed_14_0_3692 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3691_inst_req_0;
      EQ_u2_u1_3691_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3691_inst_req_1;
      EQ_u2_u1_3691_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_16_gI: SplitGuardInterface generic map(name => "ApIntEq_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : EQ_u2_u1_3702_inst 
    ApIntEq_group_17: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3680;
      EQ_u2_u1_3567_3567_delayed_14_0_3703 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3702_inst_req_0;
      EQ_u2_u1_3702_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3702_inst_req_1;
      EQ_u2_u1_3702_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_17_gI: SplitGuardInterface generic map(name => "ApIntEq_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : EQ_u2_u1_3716_inst 
    ApIntEq_group_18: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3680;
      EQ_u2_u1_3575_3575_delayed_14_0_3717 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3716_inst_req_0;
      EQ_u2_u1_3716_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3716_inst_req_1;
      EQ_u2_u1_3716_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_18_gI: SplitGuardInterface generic map(name => "ApIntEq_group_18_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "10",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : EQ_u2_u1_3730_inst 
    ApIntEq_group_19: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3680;
      EQ_u2_u1_3583_3583_delayed_14_0_3731 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3730_inst_req_0;
      EQ_u2_u1_3730_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3730_inst_req_1;
      EQ_u2_u1_3730_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_19_gI: SplitGuardInterface generic map(name => "ApIntEq_group_19_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : EQ_u2_u1_3744_inst 
    ApIntEq_group_20: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3684;
      EQ_u2_u1_3591_3591_delayed_14_0_3745 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3744_inst_req_0;
      EQ_u2_u1_3744_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3744_inst_req_1;
      EQ_u2_u1_3744_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_20_gI: SplitGuardInterface generic map(name => "ApIntEq_group_20_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : EQ_u2_u1_3758_inst 
    ApIntEq_group_21: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3684;
      EQ_u2_u1_3599_3599_delayed_14_0_3759 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3758_inst_req_0;
      EQ_u2_u1_3758_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3758_inst_req_1;
      EQ_u2_u1_3758_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_21_gI: SplitGuardInterface generic map(name => "ApIntEq_group_21_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : EQ_u2_u1_3772_inst 
    ApIntEq_group_22: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3684;
      EQ_u2_u1_3607_3607_delayed_14_0_3773 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3772_inst_req_0;
      EQ_u2_u1_3772_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3772_inst_req_1;
      EQ_u2_u1_3772_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_22_gI: SplitGuardInterface generic map(name => "ApIntEq_group_22_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "10",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : EQ_u2_u1_3786_inst 
    ApIntEq_group_23: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3684;
      EQ_u2_u1_3615_3615_delayed_14_0_3787 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3786_inst_req_0;
      EQ_u2_u1_3786_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3786_inst_req_1;
      EQ_u2_u1_3786_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_23_gI: SplitGuardInterface generic map(name => "ApIntEq_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- binary operator LSHR_u32_u32_3616_inst
    process(address1_3497) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_3497, konst_3615_wire_constant, tmp_var);
      LSHR_u32_u32_3616_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3626_inst
    process(address2_3502) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_3502, konst_3625_wire_constant, tmp_var);
      LSHR_u32_u32_3626_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3492_inst
    process(chl_out_3488, cb_3485) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_out_3488, cb_3485, tmp_var);
      MUL_u16_u16_3492_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_3833_inst
    process(chl_change_3539) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", chl_change_3539, tmp_var);
      NOT_u1_u1_3833_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_3834_inst
    process(ULT_u16_u1_3831_wire, NOT_u1_u1_3833_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ULT_u16_u1_3831_wire, NOT_u1_u1_3833_wire, tmp_var);
      continue_flag_3835 <= tmp_var; --
    end process;
    -- shared split operator group (29) : SUB_u16_u16_3531_inst 
    ApIntSub_group_29: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rb_3482;
      SUB_u16_u16_3413_3413_delayed_1_0_3532 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3531_inst_req_0;
      SUB_u16_u16_3531_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3531_inst_req_1;
      SUB_u16_u16_3531_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_29_gI: SplitGuardInterface generic map(name => "ApIntSub_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : SUB_u16_u16_3826_inst 
    ApIntSub_group_30: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= chl_out_3488;
      SUB_u16_u16_3644_3644_delayed_1_0_3827 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3826_inst_req_0;
      SUB_u16_u16_3826_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3826_inst_req_1;
      SUB_u16_u16_3826_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_30_gI: SplitGuardInterface generic map(name => "ApIntSub_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- binary operator UGE_u16_u1_3537_inst
    process(row_3517, SUB_u16_u16_3413_3413_delayed_1_0_3532) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(row_3517, SUB_u16_u16_3413_3413_delayed_1_0_3532, tmp_var);
      UGE_u16_u1_3537_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_3831_inst
    process(chl_3507, SUB_u16_u16_3644_3644_delayed_1_0_3827) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(chl_3507, SUB_u16_u16_3644_3644_delayed_1_0_3827, tmp_var);
      ULT_u16_u1_3831_wire <= tmp_var; --
    end process;
    -- shared split operator group (33) : array_obj_ref_3618_index_offset 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3617_scaled;
      array_obj_ref_3618_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3618_index_offset_req_0;
      array_obj_ref_3618_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3618_index_offset_req_1;
      array_obj_ref_3618_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : array_obj_ref_3628_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3627_scaled;
      array_obj_ref_3628_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3628_index_offset_req_0;
      array_obj_ref_3628_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3628_index_offset_req_1;
      array_obj_ref_3628_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared load operator group (0) : ptr_deref_3633_load_0 ptr_deref_3637_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3633_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3637_load_0_req_0;
      ptr_deref_3633_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3637_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3633_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3637_load_0_req_1;
      ptr_deref_3633_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3637_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3633_word_address_0 & ptr_deref_3637_word_address_0;
      ptr_deref_3633_data_0 <= data_out(127 downto 64);
      ptr_deref_3637_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3814_store_0 ptr_deref_3801_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3814_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3801_store_0_req_0;
      ptr_deref_3814_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3801_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3814_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3801_store_0_req_1;
      ptr_deref_3814_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3801_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3814_word_address_0 & ptr_deref_3801_word_address_0;
      data_in <= ptr_deref_3814_data_0 & ptr_deref_3801_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_output_pipe_3487_inst RPIPE_output_pipe_3484_inst RPIPE_output_pipe_3481_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(47 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 2 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= RPIPE_output_pipe_3487_inst_req_0;
      reqL_unguarded(1) <= RPIPE_output_pipe_3484_inst_req_0;
      reqL_unguarded(0) <= RPIPE_output_pipe_3481_inst_req_0;
      RPIPE_output_pipe_3487_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_output_pipe_3484_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_output_pipe_3481_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= RPIPE_output_pipe_3487_inst_req_1;
      reqR_unguarded(1) <= RPIPE_output_pipe_3484_inst_req_1;
      reqR_unguarded(0) <= RPIPE_output_pipe_3481_inst_req_1;
      RPIPE_output_pipe_3487_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_output_pipe_3484_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_output_pipe_3481_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      chl_out_3488 <= data_out(47 downto 32);
      cb_3485 <= data_out(31 downto 16);
      rb_3482 <= data_out(15 downto 0);
      output_pipe_read_0_gI: SplitGuardInterface generic map(name => "output_pipe_read_0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_0: InputPortRevised -- 
        generic map ( name => "output_pipe_read_0", data_width => 16,  num_reqs => 3,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(1),
          oack => output_pipe_pipe_read_ack(1),
          odata => output_pipe_pipe_read_data(31 downto 16),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_output_pipe_3640_inst RPIPE_output_pipe_3643_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_output_pipe_3640_inst_req_0;
      reqL_unguarded(0) <= RPIPE_output_pipe_3643_inst_req_0;
      RPIPE_output_pipe_3640_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_output_pipe_3643_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_output_pipe_3640_inst_req_1;
      reqR_unguarded(0) <= RPIPE_output_pipe_3643_inst_req_1;
      RPIPE_output_pipe_3640_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_output_pipe_3643_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      output_data1_3641 <= data_out(31 downto 16);
      output_data2_3644 <= data_out(15 downto 0);
      output_pipe_read_1_gI: SplitGuardInterface generic map(name => "output_pipe_read_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_1: InputPortRevised -- 
        generic map ( name => "output_pipe_read_1", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(0),
          oack => output_pipe_pipe_read_ack(0),
          odata => output_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3838_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3838_inst_req_0;
      WPIPE_input_done_pipe_3838_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3838_inst_req_1;
      WPIPE_input_done_pipe_3838_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3839_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendModule_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_1875_start: Boolean;
  signal timer_CP_1875_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_828_inst_req_0 : boolean;
  signal WPIPE_timer_req_828_inst_ack_0 : boolean;
  signal WPIPE_timer_req_828_inst_req_1 : boolean;
  signal WPIPE_timer_req_828_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_833_inst_req_0 : boolean;
  signal RPIPE_timer_resp_833_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_833_inst_req_1 : boolean;
  signal RPIPE_timer_resp_833_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_1875_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1875_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_1875_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1875_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_1875: Block -- control-path 
    signal timer_CP_1875_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_1875_elements(0) <= timer_CP_1875_start;
    timer_CP_1875_symbol <= timer_CP_1875_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_831_to_assign_stmt_834/$entry
      -- CP-element group 0: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_sample_start_
      -- CP-element group 0: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_Sample/req
      -- CP-element group 0: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_sample_start_
      -- CP-element group 0: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_Sample/rr
      -- 
    req_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1875_elements(0), ack => WPIPE_timer_req_828_inst_req_0); -- 
    rr_1902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1875_elements(0), ack => RPIPE_timer_resp_833_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_sample_completed_
      -- CP-element group 1: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_update_start_
      -- CP-element group 1: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_Sample/ack
      -- CP-element group 1: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_Update/$entry
      -- CP-element group 1: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_Update/req
      -- 
    ack_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_828_inst_ack_0, ack => timer_CP_1875_elements(1)); -- 
    req_1893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1875_elements(1), ack => WPIPE_timer_req_828_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_update_completed_
      -- CP-element group 2: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_Update/$exit
      -- CP-element group 2: 	 assign_stmt_831_to_assign_stmt_834/WPIPE_timer_req_828_Update/ack
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_828_inst_ack_1, ack => timer_CP_1875_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_sample_completed_
      -- CP-element group 3: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_update_start_
      -- CP-element group 3: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_Sample/ra
      -- CP-element group 3: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_Update/$entry
      -- CP-element group 3: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_Update/cr
      -- 
    ra_1903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_833_inst_ack_0, ack => timer_CP_1875_elements(3)); -- 
    cr_1907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1875_elements(3), ack => RPIPE_timer_resp_833_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_update_completed_
      -- CP-element group 4: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_Update/$exit
      -- CP-element group 4: 	 assign_stmt_831_to_assign_stmt_834/RPIPE_timer_resp_833_Update/ca
      -- 
    ca_1908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_833_inst_ack_1, ack => timer_CP_1875_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_831_to_assign_stmt_834/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_1875_elements(2) & timer_CP_1875_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_1875_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_830_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_830_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_833_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_833_inst_req_0;
      RPIPE_timer_resp_833_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_833_inst_req_1;
      RPIPE_timer_resp_833_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_828_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_828_inst_req_0;
      WPIPE_timer_req_828_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_828_inst_req_1;
      WPIPE_timer_req_828_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_830_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_10183_start: Boolean;
  signal timerDaemon_CP_10183_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_resp_4133_inst_req_1 : boolean;
  signal nCOUNTER_4131_4122_buf_req_1 : boolean;
  signal do_while_stmt_4116_branch_ack_1 : boolean;
  signal do_while_stmt_4116_branch_ack_0 : boolean;
  signal WPIPE_timer_resp_4133_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_4133_inst_req_0 : boolean;
  signal RPIPE_timer_req_4125_inst_ack_1 : boolean;
  signal phi_stmt_4118_req_1 : boolean;
  signal RPIPE_timer_req_4125_inst_req_1 : boolean;
  signal RPIPE_timer_req_4125_inst_ack_0 : boolean;
  signal RPIPE_timer_req_4125_inst_req_0 : boolean;
  signal nCOUNTER_4131_4122_buf_ack_0 : boolean;
  signal WPIPE_timer_resp_4133_inst_ack_1 : boolean;
  signal do_while_stmt_4116_branch_req_0 : boolean;
  signal phi_stmt_4118_ack_0 : boolean;
  signal nCOUNTER_4131_4122_buf_ack_1 : boolean;
  signal nCOUNTER_4131_4122_buf_req_0 : boolean;
  signal phi_stmt_4118_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_10183_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_10183_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_10183_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_10183_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_10183: Block -- control-path 
    signal timerDaemon_CP_10183_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_10183_elements(0) <= timerDaemon_CP_10183_start;
    timerDaemon_CP_10183_symbol <= timerDaemon_CP_10183_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_4115/branch_block_stmt_4115__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_4115/do_while_stmt_4116__entry__
      -- CP-element group 0: 	 branch_block_stmt_4115/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_4115/branch_block_stmt_4115__exit__
      -- CP-element group 1: 	 branch_block_stmt_4115/$exit
      -- CP-element group 1: 	 branch_block_stmt_4115/do_while_stmt_4116__exit__
      -- CP-element group 1: 	 $exit
      -- 
    timerDaemon_CP_10183_elements(1) <= timerDaemon_CP_10183_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116__entry__
      -- CP-element group 2: 	 branch_block_stmt_4115/do_while_stmt_4116/$entry
      -- 
    timerDaemon_CP_10183_elements(2) <= timerDaemon_CP_10183_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116__exit__
      -- 
    -- Element group timerDaemon_CP_10183_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_4115/do_while_stmt_4116/loop_back
      -- 
    -- Element group timerDaemon_CP_10183_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_4115/do_while_stmt_4116/condition_done
      -- CP-element group 5: 	 branch_block_stmt_4115/do_while_stmt_4116/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_4115/do_while_stmt_4116/loop_exit/$entry
      -- 
    timerDaemon_CP_10183_elements(5) <= timerDaemon_CP_10183_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_4115/do_while_stmt_4116/loop_body_done
      -- 
    timerDaemon_CP_10183_elements(6) <= timerDaemon_CP_10183_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_10183_elements(7) <= timerDaemon_CP_10183_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_10183_elements(8) <= timerDaemon_CP_10183_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4123_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/$entry
      -- 
    -- Element group timerDaemon_CP_10183_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/condition_evaluated
      -- 
    condition_evaluated_10207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_10207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(10), ack => do_while_stmt_4116_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(40) & timerDaemon_CP_10183_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/aggregated_phi_sample_req
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(9) & timerDaemon_CP_10183_elements(15) & timerDaemon_CP_10183_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4123_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/aggregated_phi_sample_ack
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(17) & timerDaemon_CP_10183_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(32) & timerDaemon_CP_10183_elements(16);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(18) & timerDaemon_CP_10183_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(9) & timerDaemon_CP_10183_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(9) & timerDaemon_CP_10183_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_10183_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_10183_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_loopback_trigger
      -- 
    timerDaemon_CP_10183_elements(19) <= timerDaemon_CP_10183_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_loopback_sample_req
      -- 
    phi_stmt_4118_loopback_sample_req_10222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4118_loopback_sample_req_10222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(20), ack => phi_stmt_4118_req_1); -- 
    -- Element group timerDaemon_CP_10183_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_entry_trigger
      -- 
    timerDaemon_CP_10183_elements(21) <= timerDaemon_CP_10183_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_entry_sample_req
      -- 
    phi_stmt_4118_entry_sample_req_10225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4118_entry_sample_req_10225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(22), ack => phi_stmt_4118_req_0); -- 
    -- Element group timerDaemon_CP_10183_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4118_phi_mux_ack
      -- 
    phi_stmt_4118_phi_mux_ack_10228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4118_ack_0, ack => timerDaemon_CP_10183_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/type_cast_4121_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/type_cast_4121_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/type_cast_4121_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/type_cast_4121_sample_start_
      -- 
    -- Element group timerDaemon_CP_10183_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/type_cast_4121_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/type_cast_4121_update_start_
      -- 
    -- Element group timerDaemon_CP_10183_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/type_cast_4121_update_completed__ps
      -- 
    timerDaemon_CP_10183_elements(26) <= timerDaemon_CP_10183_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/type_cast_4121_update_completed_
      -- 
    -- Element group timerDaemon_CP_10183_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_10183_elements(25), ack => timerDaemon_CP_10183_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_Sample/req
      -- 
    req_10249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(28), ack => nCOUNTER_4131_4122_buf_req_0); -- 
    -- Element group timerDaemon_CP_10183_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_update_start_
      -- CP-element group 29: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_Update/req
      -- 
    req_10254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(29), ack => nCOUNTER_4131_4122_buf_req_1); -- 
    -- Element group timerDaemon_CP_10183_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_Sample/ack
      -- 
    ack_10250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_4131_4122_buf_ack_0, ack => timerDaemon_CP_10183_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/R_nCOUNTER_4122_Update/$exit
      -- 
    ack_10255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_4131_4122_buf_ack_1, ack => timerDaemon_CP_10183_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4123_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(9) & timerDaemon_CP_10183_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_Sample/$entry
      -- 
    rr_10268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(33), ack => RPIPE_timer_req_4125_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(11) & timerDaemon_CP_10183_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_update_start_
      -- CP-element group 34: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_Update/cr
      -- 
    cr_10273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(34), ack => RPIPE_timer_req_4125_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(13) & timerDaemon_CP_10183_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_Sample/$exit
      -- 
    ra_10269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_4125_inst_ack_0, ack => timerDaemon_CP_10183_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/phi_stmt_4123_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/RPIPE_timer_req_4125_update_completed_
      -- 
    ca_10274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_4125_inst_ack_1, ack => timerDaemon_CP_10183_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_Sample/$entry
      -- 
    req_10282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(37), ack => WPIPE_timer_resp_4133_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(18) & timerDaemon_CP_10183_elements(36) & timerDaemon_CP_10183_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_Update/req
      -- CP-element group 38: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_update_start_
      -- CP-element group 38: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_Sample/$exit
      -- 
    ack_10283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_4133_inst_ack_0, ack => timerDaemon_CP_10183_elements(38)); -- 
    req_10287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10183_elements(38), ack => WPIPE_timer_resp_4133_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/WPIPE_timer_resp_4133_Update/ack
      -- 
    ack_10288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_4133_inst_ack_1, ack => timerDaemon_CP_10183_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_10183_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_10183_elements(9), ack => timerDaemon_CP_10183_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_4115/do_while_stmt_4116/do_while_stmt_4116_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10183_elements(39) & timerDaemon_CP_10183_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10183_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_4115/do_while_stmt_4116/loop_exit/ack
      -- CP-element group 42: 	 branch_block_stmt_4115/do_while_stmt_4116/loop_exit/$exit
      -- 
    ack_10293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_4116_branch_ack_0, ack => timerDaemon_CP_10183_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_4115/do_while_stmt_4116/loop_taken/ack
      -- CP-element group 43: 	 branch_block_stmt_4115/do_while_stmt_4116/loop_taken/$exit
      -- 
    ack_10297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_4116_branch_ack_1, ack => timerDaemon_CP_10183_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_4115/do_while_stmt_4116/$exit
      -- 
    timerDaemon_CP_10183_elements(44) <= timerDaemon_CP_10183_elements(3);
    timerDaemon_do_while_stmt_4116_terminator_10298: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_4116_terminator_10298", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_10183_elements(6),loop_continue => timerDaemon_CP_10183_elements(43),loop_terminate => timerDaemon_CP_10183_elements(42),loop_back => timerDaemon_CP_10183_elements(4),loop_exit => timerDaemon_CP_10183_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_4118_phi_seq_10256_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_10183_elements(21);
      timerDaemon_CP_10183_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_10183_elements(24);
      timerDaemon_CP_10183_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_10183_elements(26);
      timerDaemon_CP_10183_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_10183_elements(19);
      timerDaemon_CP_10183_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_10183_elements(30);
      timerDaemon_CP_10183_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_10183_elements(31);
      timerDaemon_CP_10183_elements(20) <= phi_mux_reqs(1);
      phi_stmt_4118_phi_seq_10256 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_4118_phi_seq_10256") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_10183_elements(11), 
          phi_sample_ack => timerDaemon_CP_10183_elements(17), 
          phi_update_req => timerDaemon_CP_10183_elements(13), 
          phi_update_ack => timerDaemon_CP_10183_elements(18), 
          phi_mux_ack => timerDaemon_CP_10183_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_10208_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_10183_elements(7);
        preds(1)  <= timerDaemon_CP_10183_elements(8);
        entry_tmerge_10208 : transition_merge -- 
          generic map(name => " entry_tmerge_10208")
          port map (preds => preds, symbol_out => timerDaemon_CP_10183_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_4118 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_4125_wire : std_logic_vector(0 downto 0);
    signal konst_4129_wire_constant : std_logic_vector(63 downto 0);
    signal konst_4137_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_4131 : std_logic_vector(63 downto 0);
    signal nCOUNTER_4131_4122_buffered : std_logic_vector(63 downto 0);
    signal req_4123 : std_logic_vector(0 downto 0);
    signal type_cast_4121_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_4129_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_4137_wire_constant <= "1";
    type_cast_4121_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_4118: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4121_wire_constant & nCOUNTER_4131_4122_buffered;
      req <= phi_stmt_4118_req_0 & phi_stmt_4118_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4118",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4118_ack_0,
          idata => idata,
          odata => COUNTER_4118,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4118
    nCOUNTER_4131_4122_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_4131_4122_buf_req_0;
      nCOUNTER_4131_4122_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_4131_4122_buf_req_1;
      nCOUNTER_4131_4122_buf_ack_1<= rack(0);
      nCOUNTER_4131_4122_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_4131_4122_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_4131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_4131_4122_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_4123
    process(RPIPE_timer_req_4125_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_4125_wire(0 downto 0);
      req_4123 <= tmp_var; -- 
    end process;
    do_while_stmt_4116_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_4137_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_4116_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_4116_branch_req_0,
          ack0 => do_while_stmt_4116_branch_ack_0,
          ack1 => do_while_stmt_4116_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_4130_inst
    process(COUNTER_4118) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_4118, konst_4129_wire_constant, tmp_var);
      nCOUNTER_4131 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_4125_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_4125_inst_req_0;
      RPIPE_timer_req_4125_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_4125_inst_req_1;
      RPIPE_timer_req_4125_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_4125_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_4133_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_4133_inst_req_0;
      WPIPE_timer_resp_4133_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_4133_inst_req_1;
      WPIPE_timer_resp_4133_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_4123(0);
      data_in <= COUNTER_4118;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(27 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(37 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(127 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_row_in :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(47 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(47 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(47 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(63 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe4_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_num_chl :  std_logic_vector(15 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(79 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(79 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(63 downto 0);
  signal sendB_in_args    : std_logic_vector(63 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(63 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendModule
  component sendModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
      output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendModule
  signal sendModule_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendModule_tag_out   : std_logic_vector(1 downto 0);
  signal sendModule_start_req : std_logic;
  signal sendModule_start_ack : std_logic;
  signal sendModule_fin_req   : std_logic;
  signal sendModule_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe2
  signal input_pipe2_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe2
  signal input_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe3
  signal input_pipe3_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe3
  signal input_pipe3_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe4
  signal input_pipe4_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe4_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe4
  signal input_pipe4_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe4_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe2
  signal kernel_pipe2_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe2
  signal kernel_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe3
  signal kernel_pipe3_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe3
  signal kernel_pipe3_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe output_pipe
  signal output_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe output_pipe
  signal output_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_row_in <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 48,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      row_in => access_T_row_in,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(19 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(2 downto 0),
      input_pipe2_pipe_write_req => input_pipe2_pipe_write_req(0 downto 0),
      input_pipe2_pipe_write_ack => input_pipe2_pipe_write_ack(0 downto 0),
      input_pipe2_pipe_write_data => input_pipe2_pipe_write_data(15 downto 0),
      input_pipe3_pipe_write_req => input_pipe3_pipe_write_req(0 downto 0),
      input_pipe3_pipe_write_ack => input_pipe3_pipe_write_ack(0 downto 0),
      input_pipe3_pipe_write_data => input_pipe3_pipe_write_data(15 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      input_pipe4_pipe_write_req => input_pipe4_pipe_write_req(0 downto 0),
      input_pipe4_pipe_write_ack => input_pipe4_pipe_write_ack(0 downto 0),
      input_pipe4_pipe_write_data => input_pipe4_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(19 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(7 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(1 downto 1),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(1 downto 1),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(31 downto 16),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(47 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(79 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(63 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe2_pipe_read_req => input_pipe2_pipe_read_req(0 downto 0),
      input_pipe2_pipe_read_ack => input_pipe2_pipe_read_ack(0 downto 0),
      input_pipe2_pipe_read_data => input_pipe2_pipe_read_data(15 downto 0),
      input_pipe3_pipe_read_req => input_pipe3_pipe_read_req(0 downto 0),
      input_pipe3_pipe_read_ack => input_pipe3_pipe_read_ack(0 downto 0),
      input_pipe3_pipe_read_data => input_pipe3_pipe_read_data(15 downto 0),
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      kernel_pipe2_pipe_read_req => kernel_pipe2_pipe_read_req(0 downto 0),
      kernel_pipe2_pipe_read_ack => kernel_pipe2_pipe_read_ack(0 downto 0),
      kernel_pipe2_pipe_read_data => kernel_pipe2_pipe_read_data(15 downto 0),
      kernel_pipe3_pipe_read_req => kernel_pipe3_pipe_read_req(0 downto 0),
      kernel_pipe3_pipe_read_ack => kernel_pipe3_pipe_read_ack(0 downto 0),
      kernel_pipe3_pipe_read_data => kernel_pipe3_pipe_read_data(15 downto 0),
      input_pipe4_pipe_read_req => input_pipe4_pipe_read_req(0 downto 0),
      input_pipe4_pipe_read_ack => input_pipe4_pipe_read_ack(0 downto 0),
      input_pipe4_pipe_read_data => input_pipe4_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(1 downto 1),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(1 downto 1),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(15 downto 8),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(0 downto 0),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(0 downto 0),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(79 downto 16);
  loadKernelChannel_num_chl <= loadKernelChannel_in_args(15 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 80,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      num_chl => loadKernelChannel_num_chl,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(1 downto 1),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(1 downto 1),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(15 downto 8),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(0 downto 0),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(0 downto 0),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(15 downto 0),
      kernel_pipe3_pipe_write_req => kernel_pipe3_pipe_write_req(0 downto 0),
      kernel_pipe3_pipe_write_ack => kernel_pipe3_pipe_write_ack(0 downto 0),
      kernel_pipe3_pipe_write_data => kernel_pipe3_pipe_write_data(15 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(15 downto 0),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(63 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(37 downto 19),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module sendModule
  sendModule_instance:sendModule-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendModule_start_req,
      start_ack => sendModule_start_ack,
      fin_req => sendModule_fin_req,
      fin_ack => sendModule_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      output_pipe_pipe_read_req => output_pipe_pipe_read_req(1 downto 0),
      output_pipe_pipe_read_ack => output_pipe_pipe_read_ack(1 downto 0),
      output_pipe_pipe_read_data => output_pipe_pipe_read_data(31 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(7 downto 0),
      tag_in => sendModule_tag_in,
      tag_out => sendModule_tag_out-- 
    ); -- 
  -- module will be run forever 
  sendModule_tag_in <= (others => '0');
  sendModule_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => sendModule_start_req, start_ack => sendModule_start_ack,  fin_req => sendModule_fin_req,  fin_ack => sendModule_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe2_pipe_read_req,
      read_ack => input_pipe2_pipe_read_ack,
      read_data => input_pipe2_pipe_read_data,
      write_req => input_pipe2_pipe_write_req,
      write_ack => input_pipe2_pipe_write_ack,
      write_data => input_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe3_pipe_read_req,
      read_ack => input_pipe3_pipe_read_ack,
      read_data => input_pipe3_pipe_read_data,
      write_req => input_pipe3_pipe_write_req,
      write_ack => input_pipe3_pipe_write_ack,
      write_data => input_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe4",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe4_pipe_read_req,
      read_ack => input_pipe4_pipe_read_ack,
      read_data => input_pipe4_pipe_read_data,
      write_req => input_pipe4_pipe_write_req,
      write_ack => input_pipe4_pipe_write_ack,
      write_data => input_pipe4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe2_pipe_read_req,
      read_ack => kernel_pipe2_pipe_read_ack,
      read_data => kernel_pipe2_pipe_read_data,
      write_req => kernel_pipe2_pipe_write_req,
      write_ack => kernel_pipe2_pipe_write_ack,
      write_data => kernel_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe3_pipe_read_req,
      read_ack => kernel_pipe3_pipe_read_ack,
      read_data => kernel_pipe3_pipe_read_data,
      write_req => kernel_pipe3_pipe_write_req,
      write_ack => kernel_pipe3_pipe_write_ack,
      write_data => kernel_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe output_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 10 --
    )
    port map( -- 
      read_req => output_pipe_pipe_read_req,
      read_ack => output_pipe_pipe_read_ack,
      read_data => output_pipe_pipe_read_data,
      write_req => output_pipe_pipe_write_req,
      write_ack => output_pipe_pipe_write_ack,
      write_data => output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 11 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
