-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_3949_start: Boolean;
  signal convTranspose_CP_3949_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1339_call_req_1 : boolean;
  signal call_stmt_1339_call_ack_1 : boolean;
  signal type_cast_1347_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1352_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1352_inst_req_1 : boolean;
  signal call_stmt_1339_call_ack_0 : boolean;
  signal call_stmt_1339_call_req_0 : boolean;
  signal RPIPE_Block1_done_1365_inst_ack_0 : boolean;
  signal type_cast_1347_inst_req_1 : boolean;
  signal type_cast_1347_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1349_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1349_inst_req_1 : boolean;
  signal call_stmt_1342_call_ack_1 : boolean;
  signal call_stmt_1342_call_req_1 : boolean;
  signal RPIPE_Block0_done_1362_inst_req_1 : boolean;
  signal call_stmt_1342_call_ack_0 : boolean;
  signal WPIPE_Block2_start_1355_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1358_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1358_inst_req_1 : boolean;
  signal call_stmt_1342_call_req_0 : boolean;
  signal WPIPE_Block2_start_1355_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1358_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1362_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1358_inst_req_0 : boolean;
  signal type_cast_1347_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1362_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1349_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1349_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1352_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1355_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1352_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1362_inst_ack_1 : boolean;
  signal call_stmt_1375_call_req_0 : boolean;
  signal call_stmt_1375_call_ack_0 : boolean;
  signal type_cast_1379_inst_req_0 : boolean;
  signal type_cast_1379_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1371_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1371_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1371_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1368_inst_ack_1 : boolean;
  signal call_stmt_1375_call_ack_1 : boolean;
  signal RPIPE_Block2_done_1368_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1365_inst_req_0 : boolean;
  signal call_stmt_1375_call_req_1 : boolean;
  signal RPIPE_Block1_done_1365_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1365_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1371_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1368_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1368_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1355_inst_req_0 : boolean;
  signal type_cast_1379_inst_req_1 : boolean;
  signal type_cast_1379_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1386_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1386_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1386_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1386_inst_ack_1 : boolean;
  signal call_stmt_1389_call_req_0 : boolean;
  signal call_stmt_1389_call_ack_0 : boolean;
  signal call_stmt_1389_call_req_1 : boolean;
  signal call_stmt_1389_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_3949_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3949_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_3949_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3949_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_3949: Block -- control-path 
    signal convTranspose_CP_3949_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    convTranspose_CP_3949_elements(0) <= convTranspose_CP_3949_start;
    convTranspose_CP_3949_symbol <= convTranspose_CP_3949_elements(32);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1337/call_stmt_1339__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1337/call_stmt_1339/$entry
      -- CP-element group 0: 	 branch_block_stmt_1337/branch_block_stmt_1337__entry__
      -- CP-element group 0: 	 branch_block_stmt_1337/$entry
      -- 
    ccr_3980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(0), ack => call_stmt_1339_call_req_1); -- 
    crr_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(0), ack => call_stmt_1339_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_sample_completed_
      -- 
    cra_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1339_call_ack_0, ack => convTranspose_CP_3949_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	19 
    -- CP-element group 2:  members (40) 
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1339__exit__
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1339/call_stmt_1339_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1339/$exit
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_Update/ccr
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_Sample/crr
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372__entry__
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_Sample/req
      -- 
    cca_3981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1339_call_ack_1, ack => convTranspose_CP_3949_elements(2)); -- 
    cr_4011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => type_cast_1347_inst_req_1); -- 
    ccr_3997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => call_stmt_1342_call_req_1); -- 
    crr_3992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => call_stmt_1342_call_req_0); -- 
    req_4062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => WPIPE_Block3_start_1358_inst_req_0); -- 
    rr_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => RPIPE_Block0_done_1362_inst_req_0); -- 
    req_4020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => WPIPE_Block0_start_1349_inst_req_0); -- 
    req_4034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => WPIPE_Block1_start_1352_inst_req_0); -- 
    rr_4104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => RPIPE_Block2_done_1368_inst_req_0); -- 
    rr_4090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => RPIPE_Block1_done_1365_inst_req_0); -- 
    rr_4118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => RPIPE_Block3_done_1371_inst_req_0); -- 
    req_4048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(2), ack => WPIPE_Block2_start_1355_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_Sample/cra
      -- CP-element group 3: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_Sample/$exit
      -- 
    cra_3993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1342_call_ack_0, ack => convTranspose_CP_3949_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/call_stmt_1342_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_Sample/$entry
      -- 
    cca_3998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1342_call_ack_1, ack => convTranspose_CP_3949_elements(4)); -- 
    rr_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(4), ack => type_cast_1347_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_Sample/$exit
      -- 
    ra_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1347_inst_ack_0, ack => convTranspose_CP_3949_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/type_cast_1347_update_completed_
      -- 
    ca_4012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1347_inst_ack_1, ack => convTranspose_CP_3949_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_Update/req
      -- CP-element group 7: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_update_start_
      -- 
    ack_4021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1349_inst_ack_0, ack => convTranspose_CP_3949_elements(7)); -- 
    req_4025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(7), ack => WPIPE_Block0_start_1349_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_Update/ack
      -- CP-element group 8: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block0_start_1349_update_completed_
      -- 
    ack_4026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1349_inst_ack_1, ack => convTranspose_CP_3949_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_Update/req
      -- CP-element group 9: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_Sample/$exit
      -- 
    ack_4035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1352_inst_ack_0, ack => convTranspose_CP_3949_elements(9)); -- 
    req_4039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(9), ack => WPIPE_Block1_start_1352_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	23 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_Update/ack
      -- CP-element group 10: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block1_start_1352_Update/$exit
      -- 
    ack_4040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1352_inst_ack_1, ack => convTranspose_CP_3949_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_Update/req
      -- CP-element group 11: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_Sample/ack
      -- CP-element group 11: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_Sample/$exit
      -- 
    ack_4049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1355_inst_ack_0, ack => convTranspose_CP_3949_elements(11)); -- 
    req_4053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(11), ack => WPIPE_Block2_start_1355_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	23 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_Update/ack
      -- CP-element group 12: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block2_start_1355_Update/$exit
      -- 
    ack_4054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1355_inst_ack_1, ack => convTranspose_CP_3949_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_Update/req
      -- CP-element group 13: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_Sample/ack
      -- CP-element group 13: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_Sample/$exit
      -- 
    ack_4063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1358_inst_ack_0, ack => convTranspose_CP_3949_elements(13)); -- 
    req_4067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(13), ack => WPIPE_Block3_start_1358_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	23 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_Update/ack
      -- CP-element group 14: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/WPIPE_Block3_start_1358_update_completed_
      -- 
    ack_4068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1358_inst_ack_1, ack => convTranspose_CP_3949_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_Update/$entry
      -- 
    ra_4077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1362_inst_ack_0, ack => convTranspose_CP_3949_elements(15)); -- 
    cr_4081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(15), ack => RPIPE_Block0_done_1362_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	23 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block0_done_1362_Update/ca
      -- 
    ca_4082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1362_inst_ack_1, ack => convTranspose_CP_3949_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_sample_completed_
      -- 
    ra_4091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1365_inst_ack_0, ack => convTranspose_CP_3949_elements(17)); -- 
    cr_4095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(17), ack => RPIPE_Block1_done_1365_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	23 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block1_done_1365_update_completed_
      -- 
    ca_4096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1365_inst_ack_1, ack => convTranspose_CP_3949_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_Update/cr
      -- 
    ra_4105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1368_inst_ack_0, ack => convTranspose_CP_3949_elements(19)); -- 
    cr_4109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(19), ack => RPIPE_Block2_done_1368_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	23 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block2_done_1368_Update/$exit
      -- 
    ca_4110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1368_inst_ack_1, ack => convTranspose_CP_3949_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_Sample/ra
      -- 
    ra_4119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1371_inst_ack_0, ack => convTranspose_CP_3949_elements(21)); -- 
    cr_4123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(21), ack => RPIPE_Block3_done_1371_inst_req_1); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/RPIPE_Block3_done_1371_update_completed_
      -- 
    ca_4124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1371_inst_ack_1, ack => convTranspose_CP_3949_elements(22)); -- 
    -- CP-element group 23:  join  fork  transition  place  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	12 
    -- CP-element group 23: 	16 
    -- CP-element group 23: 	14 
    -- CP-element group 23: 	10 
    -- CP-element group 23: 	6 
    -- CP-element group 23: 	18 
    -- CP-element group 23: 	20 
    -- CP-element group 23: 	8 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	31 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (19) 
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372/$exit
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389__entry__
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1342_to_assign_stmt_1372__exit__
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_Sample/crr
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/$entry
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_Update/ccr
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_Update/cr
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_Sample/crr
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_Update/ccr
      -- 
    crr_4135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(23), ack => call_stmt_1375_call_req_0); -- 
    ccr_4140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(23), ack => call_stmt_1375_call_req_1); -- 
    cr_4154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(23), ack => type_cast_1379_inst_req_1); -- 
    crr_4177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(23), ack => call_stmt_1389_call_req_0); -- 
    ccr_4182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(23), ack => call_stmt_1389_call_req_1); -- 
    convTranspose_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_3949_elements(12) & convTranspose_CP_3949_elements(16) & convTranspose_CP_3949_elements(14) & convTranspose_CP_3949_elements(10) & convTranspose_CP_3949_elements(6) & convTranspose_CP_3949_elements(18) & convTranspose_CP_3949_elements(20) & convTranspose_CP_3949_elements(8) & convTranspose_CP_3949_elements(22);
      gj_convTranspose_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3949_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_Sample/cra
      -- CP-element group 24: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_sample_completed_
      -- 
    cra_4136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1375_call_ack_0, ack => convTranspose_CP_3949_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_Update/cca
      -- CP-element group 25: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1375_Update/$exit
      -- 
    cca_4141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1375_call_ack_1, ack => convTranspose_CP_3949_elements(25)); -- 
    rr_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(25), ack => type_cast_1379_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_Sample/$exit
      -- 
    ra_4150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1379_inst_ack_0, ack => convTranspose_CP_3949_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/type_cast_1379_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_Sample/req
      -- 
    ca_4155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1379_inst_ack_1, ack => convTranspose_CP_3949_elements(27)); -- 
    req_4163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(27), ack => WPIPE_elapsed_time_pipe_1386_inst_req_0); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_Update/req
      -- 
    ack_4164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1386_inst_ack_0, ack => convTranspose_CP_3949_elements(28)); -- 
    req_4168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3949_elements(28), ack => WPIPE_elapsed_time_pipe_1386_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/WPIPE_elapsed_time_pipe_1386_Update/ack
      -- 
    ack_4169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1386_inst_ack_1, ack => convTranspose_CP_3949_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_Sample/cra
      -- 
    cra_4178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1389_call_ack_0, ack => convTranspose_CP_3949_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	23 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/call_stmt_1389_Update/cca
      -- 
    cca_4183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1389_call_ack_1, ack => convTranspose_CP_3949_elements(31)); -- 
    -- CP-element group 32:  join  transition  place  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: 	29 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (13) 
      -- CP-element group 32: 	 $exit
      -- CP-element group 32: 	 branch_block_stmt_1337/branch_block_stmt_1337__exit__
      -- CP-element group 32: 	 branch_block_stmt_1337/merge_stmt_1391__exit__
      -- CP-element group 32: 	 branch_block_stmt_1337/return__
      -- CP-element group 32: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389__exit__
      -- CP-element group 32: 	 branch_block_stmt_1337/$exit
      -- CP-element group 32: 	 branch_block_stmt_1337/call_stmt_1375_to_call_stmt_1389/$exit
      -- CP-element group 32: 	 branch_block_stmt_1337/return___PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_1337/return___PhiReq/$exit
      -- CP-element group 32: 	 branch_block_stmt_1337/merge_stmt_1391_PhiReqMerge
      -- CP-element group 32: 	 branch_block_stmt_1337/merge_stmt_1391_PhiAck/$entry
      -- CP-element group 32: 	 branch_block_stmt_1337/merge_stmt_1391_PhiAck/$exit
      -- CP-element group 32: 	 branch_block_stmt_1337/merge_stmt_1391_PhiAck/dummy
      -- 
    convTranspose_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_3949_elements(31) & convTranspose_CP_3949_elements(29);
      gj_convTranspose_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3949_elements(32), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call10_1369 : std_logic_vector(15 downto 0);
    signal call12_1372 : std_logic_vector(15 downto 0);
    signal call14_1375 : std_logic_vector(63 downto 0);
    signal call1_1342 : std_logic_vector(63 downto 0);
    signal call6_1363 : std_logic_vector(15 downto 0);
    signal call8_1366 : std_logic_vector(15 downto 0);
    signal call_1339 : std_logic_vector(15 downto 0);
    signal conv15_1380 : std_logic_vector(63 downto 0);
    signal conv_1348 : std_logic_vector(63 downto 0);
    signal sub_1385 : std_logic_vector(63 downto 0);
    signal type_cast_1346_wire : std_logic_vector(63 downto 0);
    signal type_cast_1378_wire : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    type_cast_1347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1347_inst_req_0;
      type_cast_1347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1347_inst_req_1;
      type_cast_1347_inst_ack_1<= rack(0);
      type_cast_1347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1346_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1348,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1379_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1379_inst_req_0;
      type_cast_1379_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1379_inst_req_1;
      type_cast_1379_inst_ack_1<= rack(0);
      type_cast_1379_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1379_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1378_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_1380,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator SUB_u64_u64_1384_inst
    process(conv15_1380, conv_1348) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv15_1380, conv_1348, tmp_var);
      sub_1385 <= tmp_var; --
    end process;
    -- unary operator type_cast_1346_inst
    process(call1_1342) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call1_1342, tmp_var);
      type_cast_1346_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1378_inst
    process(call14_1375) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call14_1375, tmp_var);
      type_cast_1378_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_Block0_done_1362_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1362_inst_req_0;
      RPIPE_Block0_done_1362_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1362_inst_req_1;
      RPIPE_Block0_done_1362_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call6_1363 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1365_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1365_inst_req_0;
      RPIPE_Block1_done_1365_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1365_inst_req_1;
      RPIPE_Block1_done_1365_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call8_1366 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1368_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1368_inst_req_0;
      RPIPE_Block2_done_1368_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1368_inst_req_1;
      RPIPE_Block2_done_1368_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call10_1369 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1371_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1371_inst_req_0;
      RPIPE_Block3_done_1371_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1371_inst_req_1;
      RPIPE_Block3_done_1371_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call12_1372 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_start_1349_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_start_1349_inst_req_0;
      WPIPE_Block0_start_1349_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_start_1349_inst_req_1;
      WPIPE_Block0_start_1349_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1339;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1352_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_start_1352_inst_req_0;
      WPIPE_Block1_start_1352_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_start_1352_inst_req_1;
      WPIPE_Block1_start_1352_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1339;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1355_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_start_1355_inst_req_0;
      WPIPE_Block2_start_1355_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_start_1355_inst_req_1;
      WPIPE_Block2_start_1355_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1339;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1358_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_start_1358_inst_req_0;
      WPIPE_Block3_start_1358_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_start_1358_inst_req_1;
      WPIPE_Block3_start_1358_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1339;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_elapsed_time_pipe_1386_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1386_inst_req_0;
      WPIPE_elapsed_time_pipe_1386_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1386_inst_req_1;
      WPIPE_elapsed_time_pipe_1386_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1385;
      elapsed_time_pipe_write_4_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1339_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1339_call_req_0;
      call_stmt_1339_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1339_call_req_1;
      call_stmt_1339_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1339 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1342_call call_stmt_1375_call 
    timer_call_group_1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1342_call_req_0;
      reqL_unguarded(0) <= call_stmt_1375_call_req_0;
      call_stmt_1342_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1375_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1342_call_req_1;
      reqR_unguarded(0) <= call_stmt_1375_call_req_1;
      call_stmt_1342_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1375_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_1_gI: SplitGuardInterface generic map(name => "timer_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call1_1342 <= data_out(127 downto 64);
      call14_1375 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1389_call 
    sendOutput_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1389_call_req_0;
      call_stmt_1389_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1389_call_req_1;
      call_stmt_1389_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_2_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_4192_start: Boolean;
  signal convTransposeA_CP_4192_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1448_load_0_ack_0 : boolean;
  signal type_cast_1469_inst_req_1 : boolean;
  signal type_cast_1469_inst_req_0 : boolean;
  signal ptr_deref_1448_load_0_req_1 : boolean;
  signal type_cast_1469_inst_ack_0 : boolean;
  signal type_cast_1455_inst_req_0 : boolean;
  signal type_cast_1455_inst_ack_0 : boolean;
  signal ptr_deref_1465_load_0_req_1 : boolean;
  signal ptr_deref_1432_load_0_req_0 : boolean;
  signal ptr_deref_1481_load_0_ack_0 : boolean;
  signal ptr_deref_1481_load_0_req_0 : boolean;
  signal ptr_deref_1465_load_0_req_0 : boolean;
  signal ptr_deref_1432_load_0_ack_1 : boolean;
  signal ptr_deref_1448_load_0_req_0 : boolean;
  signal ptr_deref_1448_load_0_ack_1 : boolean;
  signal type_cast_1436_inst_ack_1 : boolean;
  signal type_cast_1455_inst_ack_1 : boolean;
  signal type_cast_1455_inst_req_1 : boolean;
  signal ptr_deref_1481_load_0_ack_1 : boolean;
  signal ptr_deref_1481_load_0_req_1 : boolean;
  signal LOAD_padding_1451_load_0_ack_1 : boolean;
  signal ptr_deref_1432_load_0_req_1 : boolean;
  signal ptr_deref_1493_load_0_ack_0 : boolean;
  signal ptr_deref_1493_load_0_req_0 : boolean;
  signal ptr_deref_1505_load_0_ack_1 : boolean;
  signal LOAD_padding_1451_load_0_req_1 : boolean;
  signal ptr_deref_1505_load_0_req_0 : boolean;
  signal ptr_deref_1505_load_0_ack_0 : boolean;
  signal ptr_deref_1505_load_0_req_1 : boolean;
  signal ptr_deref_1493_load_0_req_1 : boolean;
  signal ptr_deref_1493_load_0_ack_1 : boolean;
  signal type_cast_1436_inst_req_1 : boolean;
  signal type_cast_1436_inst_ack_0 : boolean;
  signal type_cast_1436_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1397_inst_req_0 : boolean;
  signal LOAD_padding_1451_load_0_ack_0 : boolean;
  signal RPIPE_Block0_start_1397_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1397_inst_req_1 : boolean;
  signal LOAD_padding_1451_load_0_req_0 : boolean;
  signal RPIPE_Block0_start_1397_inst_ack_1 : boolean;
  signal type_cast_1469_inst_ack_1 : boolean;
  signal ptr_deref_1465_load_0_ack_0 : boolean;
  signal ptr_deref_1432_load_0_ack_0 : boolean;
  signal ptr_deref_1410_load_0_req_0 : boolean;
  signal ptr_deref_1410_load_0_ack_0 : boolean;
  signal ptr_deref_1410_load_0_req_1 : boolean;
  signal ptr_deref_1410_load_0_ack_1 : boolean;
  signal ptr_deref_1422_load_0_req_0 : boolean;
  signal ptr_deref_1422_load_0_ack_0 : boolean;
  signal ptr_deref_1422_load_0_req_1 : boolean;
  signal ptr_deref_1422_load_0_ack_1 : boolean;
  signal ptr_deref_1465_load_0_ack_1 : boolean;
  signal ptr_deref_1523_load_0_req_0 : boolean;
  signal ptr_deref_1523_load_0_ack_0 : boolean;
  signal ptr_deref_1523_load_0_req_1 : boolean;
  signal ptr_deref_1523_load_0_ack_1 : boolean;
  signal type_cast_1552_inst_req_0 : boolean;
  signal type_cast_1552_inst_ack_0 : boolean;
  signal type_cast_1552_inst_req_1 : boolean;
  signal type_cast_1552_inst_ack_1 : boolean;
  signal type_cast_1557_inst_req_0 : boolean;
  signal type_cast_1557_inst_ack_0 : boolean;
  signal type_cast_1557_inst_req_1 : boolean;
  signal type_cast_1557_inst_ack_1 : boolean;
  signal type_cast_1679_inst_req_0 : boolean;
  signal type_cast_1679_inst_ack_0 : boolean;
  signal type_cast_1679_inst_req_1 : boolean;
  signal type_cast_1679_inst_ack_1 : boolean;
  signal type_cast_1709_inst_req_0 : boolean;
  signal type_cast_1709_inst_ack_0 : boolean;
  signal type_cast_1709_inst_req_1 : boolean;
  signal type_cast_1709_inst_ack_1 : boolean;
  signal array_obj_ref_1715_index_offset_req_0 : boolean;
  signal array_obj_ref_1715_index_offset_ack_0 : boolean;
  signal array_obj_ref_1715_index_offset_req_1 : boolean;
  signal array_obj_ref_1715_index_offset_ack_1 : boolean;
  signal addr_of_1716_final_reg_req_0 : boolean;
  signal addr_of_1716_final_reg_ack_0 : boolean;
  signal addr_of_1716_final_reg_req_1 : boolean;
  signal addr_of_1716_final_reg_ack_1 : boolean;
  signal ptr_deref_1720_load_0_req_0 : boolean;
  signal ptr_deref_1720_load_0_ack_0 : boolean;
  signal ptr_deref_1720_load_0_req_1 : boolean;
  signal ptr_deref_1720_load_0_ack_1 : boolean;
  signal type_cast_1740_inst_req_0 : boolean;
  signal type_cast_1740_inst_ack_0 : boolean;
  signal type_cast_1740_inst_req_1 : boolean;
  signal type_cast_1740_inst_ack_1 : boolean;
  signal array_obj_ref_1746_index_offset_req_0 : boolean;
  signal array_obj_ref_1746_index_offset_ack_0 : boolean;
  signal array_obj_ref_1746_index_offset_req_1 : boolean;
  signal array_obj_ref_1746_index_offset_ack_1 : boolean;
  signal addr_of_1747_final_reg_req_0 : boolean;
  signal addr_of_1747_final_reg_ack_0 : boolean;
  signal addr_of_1747_final_reg_req_1 : boolean;
  signal addr_of_1747_final_reg_ack_1 : boolean;
  signal ptr_deref_1750_store_0_req_0 : boolean;
  signal ptr_deref_1750_store_0_ack_0 : boolean;
  signal ptr_deref_1750_store_0_req_1 : boolean;
  signal ptr_deref_1750_store_0_ack_1 : boolean;
  signal type_cast_1756_inst_req_0 : boolean;
  signal type_cast_1756_inst_ack_0 : boolean;
  signal type_cast_1756_inst_req_1 : boolean;
  signal type_cast_1756_inst_ack_1 : boolean;
  signal if_stmt_1769_branch_req_0 : boolean;
  signal if_stmt_1769_branch_ack_1 : boolean;
  signal if_stmt_1769_branch_ack_0 : boolean;
  signal type_cast_1793_inst_req_0 : boolean;
  signal type_cast_1793_inst_ack_0 : boolean;
  signal type_cast_1793_inst_req_1 : boolean;
  signal type_cast_1793_inst_ack_1 : boolean;
  signal type_cast_1802_inst_req_0 : boolean;
  signal type_cast_1802_inst_ack_0 : boolean;
  signal type_cast_1802_inst_req_1 : boolean;
  signal type_cast_1802_inst_ack_1 : boolean;
  signal type_cast_1819_inst_req_0 : boolean;
  signal type_cast_1819_inst_ack_0 : boolean;
  signal type_cast_1819_inst_req_1 : boolean;
  signal type_cast_1819_inst_ack_1 : boolean;
  signal if_stmt_1826_branch_req_0 : boolean;
  signal if_stmt_1826_branch_ack_1 : boolean;
  signal if_stmt_1826_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1834_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1834_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1834_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1834_inst_ack_1 : boolean;
  signal phi_stmt_1533_req_0 : boolean;
  signal phi_stmt_1540_req_0 : boolean;
  signal type_cast_1539_inst_req_0 : boolean;
  signal type_cast_1539_inst_ack_0 : boolean;
  signal type_cast_1539_inst_req_1 : boolean;
  signal type_cast_1539_inst_ack_1 : boolean;
  signal phi_stmt_1533_req_1 : boolean;
  signal type_cast_1546_inst_req_0 : boolean;
  signal type_cast_1546_inst_ack_0 : boolean;
  signal type_cast_1546_inst_req_1 : boolean;
  signal type_cast_1546_inst_ack_1 : boolean;
  signal phi_stmt_1540_req_1 : boolean;
  signal phi_stmt_1533_ack_0 : boolean;
  signal phi_stmt_1540_ack_0 : boolean;
  signal type_cast_1669_inst_req_0 : boolean;
  signal type_cast_1669_inst_ack_0 : boolean;
  signal type_cast_1669_inst_req_1 : boolean;
  signal type_cast_1669_inst_ack_1 : boolean;
  signal phi_stmt_1663_req_1 : boolean;
  signal phi_stmt_1663_req_0 : boolean;
  signal phi_stmt_1663_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_4192_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_4192_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_4192_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_4192_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_4192: Block -- control-path 
    signal convTransposeA_CP_4192_elements: BooleanArray(88 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_4192_elements(0) <= convTransposeA_CP_4192_start;
    convTransposeA_CP_4192_symbol <= convTransposeA_CP_4192_elements(68);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1395/$entry
      -- CP-element group 0: 	 branch_block_stmt_1395/branch_block_stmt_1395__entry__
      -- CP-element group 0: 	 branch_block_stmt_1395/assign_stmt_1398__entry__
      -- CP-element group 0: 	 branch_block_stmt_1395/assign_stmt_1398/$entry
      -- CP-element group 0: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_Sample/rr
      -- 
    rr_4240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(0), ack => RPIPE_Block0_start_1397_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_Update/cr
      -- 
    ra_4241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1397_inst_ack_0, ack => convTransposeA_CP_4192_elements(1)); -- 
    cr_4245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(1), ack => RPIPE_Block0_start_1397_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1398__exit__
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530__entry__
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1398/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1398/RPIPE_Block0_start_1397_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/word_access_complete/word_0/cr
      -- 
    ca_4246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1397_inst_ack_1, ack => convTransposeA_CP_4192_elements(2)); -- 
    cr_4573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => type_cast_1469_inst_req_1); -- 
    cr_4457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1448_load_0_req_1); -- 
    cr_4554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1465_load_0_req_1); -- 
    rr_4382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1432_load_0_req_0); -- 
    rr_4607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1481_load_0_req_0); -- 
    rr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1465_load_0_req_0); -- 
    rr_4446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1448_load_0_req_0); -- 
    cr_4509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => type_cast_1455_inst_req_1); -- 
    cr_4618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1481_load_0_req_1); -- 
    cr_4393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1432_load_0_req_1); -- 
    rr_4657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1493_load_0_req_0); -- 
    cr_4490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => LOAD_padding_1451_load_0_req_1); -- 
    rr_4707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1505_load_0_req_0); -- 
    cr_4718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1505_load_0_req_1); -- 
    cr_4668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1493_load_0_req_1); -- 
    cr_4412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => type_cast_1436_inst_req_1); -- 
    rr_4479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => LOAD_padding_1451_load_0_req_0); -- 
    rr_4282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1410_load_0_req_0); -- 
    cr_4293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1410_load_0_req_1); -- 
    rr_4332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1422_load_0_req_0); -- 
    cr_4343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1422_load_0_req_1); -- 
    rr_4757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1523_load_0_req_0); -- 
    cr_4768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(2), ack => ptr_deref_1523_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Sample/word_access_start/word_0/ra
      -- 
    ra_4283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1410_load_0_ack_0, ack => convTransposeA_CP_4192_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	29 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/ptr_deref_1410_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/ptr_deref_1410_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/ptr_deref_1410_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1410_Update/ptr_deref_1410_Merge/merge_ack
      -- 
    ca_4294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1410_load_0_ack_1, ack => convTransposeA_CP_4192_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Sample/word_access_start/word_0/ra
      -- 
    ra_4333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1422_load_0_ack_0, ack => convTransposeA_CP_4192_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	29 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/ptr_deref_1422_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/ptr_deref_1422_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/ptr_deref_1422_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1422_Update/ptr_deref_1422_Merge/merge_ack
      -- 
    ca_4344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1422_load_0_ack_1, ack => convTransposeA_CP_4192_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_sample_completed_
      -- 
    ra_4383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1432_load_0_ack_0, ack => convTransposeA_CP_4192_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/ptr_deref_1432_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/ptr_deref_1432_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/ptr_deref_1432_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/ptr_deref_1432_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1432_update_completed_
      -- 
    ca_4394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1432_load_0_ack_1, ack => convTransposeA_CP_4192_elements(8)); -- 
    rr_4407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(8), ack => type_cast_1436_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_Sample/ra
      -- 
    ra_4408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1436_inst_ack_0, ack => convTransposeA_CP_4192_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1436_Update/$exit
      -- 
    ca_4413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1436_inst_ack_1, ack => convTransposeA_CP_4192_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Sample/word_access_start/word_0/ra
      -- CP-element group 11: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Sample/word_access_start/word_0/$exit
      -- 
    ra_4447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1448_load_0_ack_0, ack => convTransposeA_CP_4192_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/ptr_deref_1448_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/ptr_deref_1448_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/ptr_deref_1448_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1448_Update/ptr_deref_1448_Merge/$entry
      -- 
    ca_4458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1448_load_0_ack_1, ack => convTransposeA_CP_4192_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Sample/word_access_start/$exit
      -- 
    ra_4480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1451_load_0_ack_0, ack => convTransposeA_CP_4192_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/LOAD_padding_1451_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/LOAD_padding_1451_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/LOAD_padding_1451_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/LOAD_padding_1451_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/LOAD_padding_1451_Update/$exit
      -- 
    ca_4491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1451_load_0_ack_1, ack => convTransposeA_CP_4192_elements(14)); -- 
    rr_4504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(14), ack => type_cast_1455_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_sample_completed_
      -- 
    ra_4505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_0, ack => convTransposeA_CP_4192_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1455_Update/$exit
      -- 
    ca_4510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_1, ack => convTransposeA_CP_4192_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Sample/word_access_start/word_0/ra
      -- 
    ra_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1465_load_0_ack_0, ack => convTransposeA_CP_4192_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/ptr_deref_1465_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/ptr_deref_1465_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/ptr_deref_1465_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/ptr_deref_1465_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1465_Update/word_access_complete/word_0/ca
      -- 
    ca_4555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1465_load_0_ack_1, ack => convTransposeA_CP_4192_elements(18)); -- 
    rr_4568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(18), ack => type_cast_1469_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_sample_completed_
      -- 
    ra_4569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1469_inst_ack_0, ack => convTransposeA_CP_4192_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/type_cast_1469_Update/ca
      -- 
    ca_4574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1469_inst_ack_1, ack => convTransposeA_CP_4192_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Sample/word_access_start/word_0/ra
      -- CP-element group 21: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_sample_completed_
      -- 
    ra_4608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1481_load_0_ack_0, ack => convTransposeA_CP_4192_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/ptr_deref_1481_Merge/merge_ack
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/ptr_deref_1481_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/ptr_deref_1481_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/ptr_deref_1481_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1481_update_completed_
      -- 
    ca_4619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1481_load_0_ack_1, ack => convTransposeA_CP_4192_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Sample/word_access_start/word_0/ra
      -- CP-element group 23: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Sample/$exit
      -- 
    ra_4658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1493_load_0_ack_0, ack => convTransposeA_CP_4192_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/ptr_deref_1493_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/ptr_deref_1493_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/ptr_deref_1493_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1493_Update/ptr_deref_1493_Merge/$entry
      -- 
    ca_4669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1493_load_0_ack_1, ack => convTransposeA_CP_4192_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_sample_completed_
      -- 
    ra_4708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1505_load_0_ack_0, ack => convTransposeA_CP_4192_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/ptr_deref_1505_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/ptr_deref_1505_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/ptr_deref_1505_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1505_Update/ptr_deref_1505_Merge/merge_ack
      -- 
    ca_4719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1505_load_0_ack_1, ack => convTransposeA_CP_4192_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Sample/word_access_start/word_0/ra
      -- 
    ra_4758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1523_load_0_ack_0, ack => convTransposeA_CP_4192_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/ptr_deref_1523_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/ptr_deref_1523_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/ptr_deref_1523_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/ptr_deref_1523_Update/ptr_deref_1523_Merge/merge_ack
      -- 
    ca_4769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1523_load_0_ack_1, ack => convTransposeA_CP_4192_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	4 
    -- CP-element group 29: 	6 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	69 
    -- CP-element group 29: 	70 
    -- CP-element group 29:  members (8) 
      -- CP-element group 29: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530__exit__
      -- CP-element group 29: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_1395/assign_stmt_1407_to_assign_stmt_1530/$exit
      -- CP-element group 29: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/$entry
      -- CP-element group 29: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/$entry
      -- CP-element group 29: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/$entry
      -- 
    convTransposeA_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(4) & convTransposeA_CP_4192_elements(6) & convTransposeA_CP_4192_elements(10) & convTransposeA_CP_4192_elements(12) & convTransposeA_CP_4192_elements(16) & convTransposeA_CP_4192_elements(20) & convTransposeA_CP_4192_elements(22) & convTransposeA_CP_4192_elements(24) & convTransposeA_CP_4192_elements(26) & convTransposeA_CP_4192_elements(28);
      gj_convTransposeA_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	82 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_Sample/ra
      -- 
    ra_4786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1552_inst_ack_0, ack => convTransposeA_CP_4192_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	82 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_Update/ca
      -- 
    ca_4791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1552_inst_ack_1, ack => convTransposeA_CP_4192_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	82 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_Sample/ra
      -- 
    ra_4800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1557_inst_ack_0, ack => convTransposeA_CP_4192_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	82 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_Update/ca
      -- 
    ca_4805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1557_inst_ack_1, ack => convTransposeA_CP_4192_elements(33)); -- 
    -- CP-element group 34:  join  transition  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	86 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660__exit__
      -- CP-element group 34: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/$exit
      -- CP-element group 34: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1663/$entry
      -- CP-element group 34: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/$entry
      -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(31) & convTransposeA_CP_4192_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_Sample/ra
      -- 
    ra_4817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1679_inst_ack_0, ack => convTransposeA_CP_4192_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	88 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	45 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_Sample/rr
      -- 
    ca_4822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1679_inst_ack_1, ack => convTransposeA_CP_4192_elements(36)); -- 
    rr_4830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(36), ack => type_cast_1709_inst_req_0); -- 
    rr_4940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(36), ack => type_cast_1740_inst_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_Sample/ra
      -- 
    ra_4831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1709_inst_ack_0, ack => convTransposeA_CP_4192_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	88 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (16) 
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_resized_1
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_scaled_1
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_computed_1
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_resize_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_resize_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_resize_1/index_resize_req
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_resize_1/index_resize_ack
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_scale_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_scale_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_scale_1/scale_rename_req
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_index_scale_1/scale_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_Sample/req
      -- 
    ca_4836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1709_inst_ack_1, ack => convTransposeA_CP_4192_elements(38)); -- 
    req_4861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(38), ack => array_obj_ref_1715_index_offset_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	56 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_sample_complete
      -- CP-element group 39: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_Sample/ack
      -- 
    ack_4862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1715_index_offset_ack_0, ack => convTransposeA_CP_4192_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	88 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (11) 
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_root_address_calculated
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_offset_calculated
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_base_plus_offset/$entry
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_base_plus_offset/$exit
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_base_plus_offset/sum_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_base_plus_offset/sum_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_request/$entry
      -- CP-element group 40: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_request/req
      -- 
    ack_4867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1715_index_offset_ack_1, ack => convTransposeA_CP_4192_elements(40)); -- 
    req_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(40), ack => addr_of_1716_final_reg_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_request/$exit
      -- CP-element group 41: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_request/ack
      -- 
    ack_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1716_final_reg_ack_0, ack => convTransposeA_CP_4192_elements(41)); -- 
    -- CP-element group 42:  join  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	88 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (24) 
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_complete/$exit
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_complete/ack
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_word_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_address_resized
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_addr_resize/$entry
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_addr_resize/$exit
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_addr_resize/base_resize_req
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_addr_resize/base_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_word_addrgen/$entry
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_word_addrgen/$exit
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_word_addrgen/root_register_req
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_word_addrgen/root_register_ack
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Sample/word_access_start/word_0/rr
      -- 
    ack_4882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1716_final_reg_ack_1, ack => convTransposeA_CP_4192_elements(42)); -- 
    rr_4915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(42), ack => ptr_deref_1720_load_0_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Sample/word_access_start/word_0/ra
      -- 
    ra_4916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1720_load_0_ack_0, ack => convTransposeA_CP_4192_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	88 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	51 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/word_access_complete/word_0/ca
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/ptr_deref_1720_Merge/$entry
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/ptr_deref_1720_Merge/$exit
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/ptr_deref_1720_Merge/merge_req
      -- CP-element group 44: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/ptr_deref_1720_Merge/merge_ack
      -- 
    ca_4927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1720_load_0_ack_1, ack => convTransposeA_CP_4192_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	36 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_Sample/ra
      -- 
    ra_4941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1740_inst_ack_0, ack => convTransposeA_CP_4192_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	88 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (16) 
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_resized_1
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_scaled_1
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_computed_1
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_resize_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_resize_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_resize_1/index_resize_req
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_resize_1/index_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_scale_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_scale_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_scale_1/scale_rename_req
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_index_scale_1/scale_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_Sample/req
      -- 
    ca_4946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1740_inst_ack_1, ack => convTransposeA_CP_4192_elements(46)); -- 
    req_4971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(46), ack => array_obj_ref_1746_index_offset_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_sample_complete
      -- CP-element group 47: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_Sample/ack
      -- 
    ack_4972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1746_index_offset_ack_0, ack => convTransposeA_CP_4192_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	88 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (11) 
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_request/$entry
      -- CP-element group 48: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_request/req
      -- 
    ack_4977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1746_index_offset_ack_1, ack => convTransposeA_CP_4192_elements(48)); -- 
    req_4986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(48), ack => addr_of_1747_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_request/ack
      -- 
    ack_4987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1747_final_reg_ack_0, ack => convTransposeA_CP_4192_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	88 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_word_addrgen/root_register_ack
      -- 
    ack_4992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1747_final_reg_ack_1, ack => convTransposeA_CP_4192_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	44 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/ptr_deref_1750_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/ptr_deref_1750_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/ptr_deref_1750_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/ptr_deref_1750_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/word_access_start/word_0/rr
      -- 
    rr_5030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(51), ack => ptr_deref_1750_store_0_req_0); -- 
    convTransposeA_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(44) & convTransposeA_CP_4192_elements(50);
      gj_convTransposeA_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Sample/word_access_start/word_0/ra
      -- 
    ra_5031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1750_store_0_ack_0, ack => convTransposeA_CP_4192_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	88 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Update/word_access_complete/word_0/ca
      -- 
    ca_5042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1750_store_0_ack_1, ack => convTransposeA_CP_4192_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	88 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_Sample/ra
      -- 
    ra_5051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1756_inst_ack_0, ack => convTransposeA_CP_4192_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	88 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_Update/ca
      -- 
    ca_5056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1756_inst_ack_1, ack => convTransposeA_CP_4192_elements(55)); -- 
    -- CP-element group 56:  branch  join  transition  place  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: 	47 
    -- CP-element group 56: 	53 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (10) 
      -- CP-element group 56: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768__exit__
      -- CP-element group 56: 	 branch_block_stmt_1395/if_stmt_1769__entry__
      -- CP-element group 56: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/$exit
      -- CP-element group 56: 	 branch_block_stmt_1395/if_stmt_1769_dead_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1395/if_stmt_1769_eval_test/$entry
      -- CP-element group 56: 	 branch_block_stmt_1395/if_stmt_1769_eval_test/$exit
      -- CP-element group 56: 	 branch_block_stmt_1395/if_stmt_1769_eval_test/branch_req
      -- CP-element group 56: 	 branch_block_stmt_1395/R_cmp_1770_place
      -- CP-element group 56: 	 branch_block_stmt_1395/if_stmt_1769_if_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1395/if_stmt_1769_else_link/$entry
      -- 
    branch_req_5064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(56), ack => if_stmt_1769_branch_req_0); -- 
    convTransposeA_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(39) & convTransposeA_CP_4192_elements(47) & convTransposeA_CP_4192_elements(53) & convTransposeA_CP_4192_elements(55);
      gj_convTransposeA_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	83 
    -- CP-element group 57: 	84 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1395/merge_stmt_1775__exit__
      -- CP-element group 57: 	 branch_block_stmt_1395/assign_stmt_1781__entry__
      -- CP-element group 57: 	 branch_block_stmt_1395/assign_stmt_1781__exit__
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody
      -- CP-element group 57: 	 branch_block_stmt_1395/if_stmt_1769_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1395/if_stmt_1769_if_link/if_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1395/whilex_xbody_ifx_xthen
      -- CP-element group 57: 	 branch_block_stmt_1395/assign_stmt_1781/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/assign_stmt_1781/$exit
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1395/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1395/merge_stmt_1775_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1395/merge_stmt_1775_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1395/merge_stmt_1775_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1395/merge_stmt_1775_PhiAck/dummy
      -- 
    if_choice_transition_5069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1769_branch_ack_1, ack => convTransposeA_CP_4192_elements(57)); -- 
    rr_5252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(57), ack => type_cast_1669_inst_req_0); -- 
    cr_5257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(57), ack => type_cast_1669_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	62 
    -- CP-element group 58: 	64 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_1395/merge_stmt_1783__exit__
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825__entry__
      -- CP-element group 58: 	 branch_block_stmt_1395/if_stmt_1769_else_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1395/if_stmt_1769_else_link/else_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1395/whilex_xbody_ifx_xelse
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/$entry
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1395/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1395/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1395/merge_stmt_1783_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1395/merge_stmt_1783_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1395/merge_stmt_1783_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1395/merge_stmt_1783_PhiAck/dummy
      -- 
    else_choice_transition_5073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1769_branch_ack_0, ack => convTransposeA_CP_4192_elements(58)); -- 
    rr_5089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(58), ack => type_cast_1793_inst_req_0); -- 
    cr_5094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(58), ack => type_cast_1793_inst_req_1); -- 
    cr_5108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(58), ack => type_cast_1802_inst_req_1); -- 
    cr_5122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(58), ack => type_cast_1819_inst_req_1); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_Sample/ra
      -- 
    ra_5090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1793_inst_ack_0, ack => convTransposeA_CP_4192_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1793_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_Sample/rr
      -- 
    ca_5095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1793_inst_ack_1, ack => convTransposeA_CP_4192_elements(60)); -- 
    rr_5103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(60), ack => type_cast_1802_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_Sample/ra
      -- 
    ra_5104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_0, ack => convTransposeA_CP_4192_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	58 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1802_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_Sample/rr
      -- 
    ca_5109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_1, ack => convTransposeA_CP_4192_elements(62)); -- 
    rr_5117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(62), ack => type_cast_1819_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_Sample/ra
      -- 
    ra_5118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1819_inst_ack_0, ack => convTransposeA_CP_4192_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	58 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825__exit__
      -- CP-element group 64: 	 branch_block_stmt_1395/if_stmt_1826__entry__
      -- CP-element group 64: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/$exit
      -- CP-element group 64: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1395/assign_stmt_1789_to_assign_stmt_1825/type_cast_1819_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_1395/if_stmt_1826_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1395/if_stmt_1826_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_1395/if_stmt_1826_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_1395/if_stmt_1826_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_1395/R_cmp77_1827_place
      -- CP-element group 64: 	 branch_block_stmt_1395/if_stmt_1826_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1395/if_stmt_1826_else_link/$entry
      -- 
    ca_5123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1819_inst_ack_1, ack => convTransposeA_CP_4192_elements(64)); -- 
    branch_req_5131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(64), ack => if_stmt_1826_branch_req_0); -- 
    -- CP-element group 65:  merge  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (15) 
      -- CP-element group 65: 	 branch_block_stmt_1395/merge_stmt_1832__exit__
      -- CP-element group 65: 	 branch_block_stmt_1395/assign_stmt_1836__entry__
      -- CP-element group 65: 	 branch_block_stmt_1395/if_stmt_1826_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1395/if_stmt_1826_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1395/ifx_xelse_whilex_xend
      -- CP-element group 65: 	 branch_block_stmt_1395/assign_stmt_1836/$entry
      -- CP-element group 65: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1395/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1395/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_1395/merge_stmt_1832_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_1395/merge_stmt_1832_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_1395/merge_stmt_1832_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1395/merge_stmt_1832_PhiAck/dummy
      -- 
    if_choice_transition_5136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1826_branch_ack_1, ack => convTransposeA_CP_4192_elements(65)); -- 
    req_5153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(65), ack => WPIPE_Block0_done_1834_inst_req_0); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	72 
    -- CP-element group 66: 	73 
    -- CP-element group 66: 	75 
    -- CP-element group 66: 	76 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_1395/if_stmt_1826_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_1395/if_stmt_1826_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1826_branch_ack_0, ack => convTransposeA_CP_4192_elements(66)); -- 
    rr_5197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(66), ack => type_cast_1539_inst_req_0); -- 
    cr_5202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(66), ack => type_cast_1539_inst_req_1); -- 
    rr_5220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(66), ack => type_cast_1546_inst_req_0); -- 
    cr_5225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(66), ack => type_cast_1546_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_Update/req
      -- 
    ack_5154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1834_inst_ack_0, ack => convTransposeA_CP_4192_elements(67)); -- 
    req_5158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(67), ack => WPIPE_Block0_done_1834_inst_req_1); -- 
    -- CP-element group 68:  transition  place  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_1395/$exit
      -- CP-element group 68: 	 branch_block_stmt_1395/branch_block_stmt_1395__exit__
      -- CP-element group 68: 	 branch_block_stmt_1395/assign_stmt_1836__exit__
      -- CP-element group 68: 	 branch_block_stmt_1395/return__
      -- CP-element group 68: 	 branch_block_stmt_1395/merge_stmt_1838__exit__
      -- CP-element group 68: 	 branch_block_stmt_1395/assign_stmt_1836/$exit
      -- CP-element group 68: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1395/assign_stmt_1836/WPIPE_Block0_done_1834_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1395/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_1395/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_1395/merge_stmt_1838_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_1395/merge_stmt_1838_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_1395/merge_stmt_1838_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_1395/merge_stmt_1838_PhiAck/dummy
      -- 
    ack_5159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1834_inst_ack_1, ack => convTransposeA_CP_4192_elements(68)); -- 
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	29 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/$exit
      -- CP-element group 69: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1537_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_req
      -- 
    phi_stmt_1533_req_5170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1533_req_5170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(69), ack => phi_stmt_1533_req_0); -- 
    -- Element group convTransposeA_CP_4192_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_4192_elements(29), ack => convTransposeA_CP_4192_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  transition  output  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/$exit
      -- CP-element group 70: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1544_konst_delay_trans
      -- CP-element group 70: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_req
      -- 
    phi_stmt_1540_req_5178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1540_req_5178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(70), ack => phi_stmt_1540_req_0); -- 
    -- Element group convTransposeA_CP_4192_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convTransposeA_CP_4192_elements(29), ack => convTransposeA_CP_4192_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	79 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1395/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(69) & convTransposeA_CP_4192_elements(70);
      gj_convTransposeA_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	66 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/Sample/ra
      -- 
    ra_5198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1539_inst_ack_0, ack => convTransposeA_CP_4192_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/Update/ca
      -- 
    ca_5203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1539_inst_ack_1, ack => convTransposeA_CP_4192_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	78 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/$exit
      -- CP-element group 74: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/$exit
      -- CP-element group 74: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1539/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1533/phi_stmt_1533_req
      -- 
    phi_stmt_1533_req_5204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1533_req_5204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(74), ack => phi_stmt_1533_req_1); -- 
    convTransposeA_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(72) & convTransposeA_CP_4192_elements(73);
      gj_convTransposeA_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	66 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/Sample/ra
      -- 
    ra_5221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1546_inst_ack_0, ack => convTransposeA_CP_4192_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	66 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/Update/ca
      -- 
    ca_5226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1546_inst_ack_1, ack => convTransposeA_CP_4192_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/$exit
      -- CP-element group 77: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/$exit
      -- CP-element group 77: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_sources/type_cast_1546/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1540/phi_stmt_1540_req
      -- 
    phi_stmt_1540_req_5227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1540_req_5227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(77), ack => phi_stmt_1540_req_1); -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(75) & convTransposeA_CP_4192_elements(76);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	74 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1395/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(74) & convTransposeA_CP_4192_elements(77);
      gj_convTransposeA_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  merge  fork  transition  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	71 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1395/merge_stmt_1532_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_1395/merge_stmt_1532_PhiAck/$entry
      -- 
    convTransposeA_CP_4192_elements(79) <= OrReduce(convTransposeA_CP_4192_elements(71) & convTransposeA_CP_4192_elements(78));
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1395/merge_stmt_1532_PhiAck/phi_stmt_1533_ack
      -- 
    phi_stmt_1533_ack_5232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1533_ack_0, ack => convTransposeA_CP_4192_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1395/merge_stmt_1532_PhiAck/phi_stmt_1540_ack
      -- 
    phi_stmt_1540_ack_5233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1540_ack_0, ack => convTransposeA_CP_4192_elements(81)); -- 
    -- CP-element group 82:  join  fork  transition  place  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	30 
    -- CP-element group 82: 	31 
    -- CP-element group 82: 	32 
    -- CP-element group 82: 	33 
    -- CP-element group 82:  members (16) 
      -- CP-element group 82: 	 branch_block_stmt_1395/merge_stmt_1532__exit__
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660__entry__
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/$entry
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1552_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1395/assign_stmt_1553_to_assign_stmt_1660/type_cast_1557_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1395/merge_stmt_1532_PhiAck/$exit
      -- 
    rr_4785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(82), ack => type_cast_1552_inst_req_0); -- 
    cr_4790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(82), ack => type_cast_1552_inst_req_1); -- 
    rr_4799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(82), ack => type_cast_1557_inst_req_0); -- 
    cr_4804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(82), ack => type_cast_1557_inst_req_1); -- 
    convTransposeA_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(80) & convTransposeA_CP_4192_elements(81);
      gj_convTransposeA_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	57 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/Sample/ra
      -- 
    ra_5253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1669_inst_ack_0, ack => convTransposeA_CP_4192_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	57 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/Update/ca
      -- 
    ca_5258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1669_inst_ack_1, ack => convTransposeA_CP_4192_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/$exit
      -- CP-element group 85: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/$exit
      -- CP-element group 85: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1669/SplitProtocol/$exit
      -- CP-element group 85: 	 branch_block_stmt_1395/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_req
      -- 
    phi_stmt_1663_req_5259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1663_req_5259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(85), ack => phi_stmt_1663_req_1); -- 
    convTransposeA_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4192_elements(83) & convTransposeA_CP_4192_elements(84);
      gj_convTransposeA_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4192_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  output  delay-element  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	34 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1663/$exit
      -- CP-element group 86: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_sources/type_cast_1667_konst_delay_trans
      -- CP-element group 86: 	 branch_block_stmt_1395/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1663/phi_stmt_1663_req
      -- 
    phi_stmt_1663_req_5270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1663_req_5270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(86), ack => phi_stmt_1663_req_0); -- 
    -- Element group convTransposeA_CP_4192_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => convTransposeA_CP_4192_elements(34), ack => convTransposeA_CP_4192_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  merge  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1395/merge_stmt_1662_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_1395/merge_stmt_1662_PhiAck/$entry
      -- 
    convTransposeA_CP_4192_elements(87) <= OrReduce(convTransposeA_CP_4192_elements(85) & convTransposeA_CP_4192_elements(86));
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	36 
    -- CP-element group 88: 	38 
    -- CP-element group 88: 	40 
    -- CP-element group 88: 	42 
    -- CP-element group 88: 	44 
    -- CP-element group 88: 	46 
    -- CP-element group 88: 	48 
    -- CP-element group 88: 	50 
    -- CP-element group 88: 	53 
    -- CP-element group 88: 	54 
    -- CP-element group 88: 	55 
    -- CP-element group 88:  members (45) 
      -- CP-element group 88: 	 branch_block_stmt_1395/merge_stmt_1662__exit__
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768__entry__
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1679_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1709_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1715_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1716_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1720_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1740_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/array_obj_ref_1746_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/addr_of_1747_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/ptr_deref_1750_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1395/assign_stmt_1676_to_assign_stmt_1768/type_cast_1756_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1395/merge_stmt_1662_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1395/merge_stmt_1662_PhiAck/phi_stmt_1663_ack
      -- 
    phi_stmt_1663_ack_5275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1663_ack_0, ack => convTransposeA_CP_4192_elements(88)); -- 
    rr_4816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => type_cast_1679_inst_req_0); -- 
    cr_4821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => type_cast_1679_inst_req_1); -- 
    cr_4835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => type_cast_1709_inst_req_1); -- 
    req_4866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => array_obj_ref_1715_index_offset_req_1); -- 
    req_4881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => addr_of_1716_final_reg_req_1); -- 
    cr_4926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => ptr_deref_1720_load_0_req_1); -- 
    cr_4945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => type_cast_1740_inst_req_1); -- 
    req_4976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => array_obj_ref_1746_index_offset_req_1); -- 
    req_4991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => addr_of_1747_final_reg_req_1); -- 
    cr_5041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => ptr_deref_1750_store_0_req_1); -- 
    rr_5050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => type_cast_1756_inst_req_0); -- 
    cr_5055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4192_elements(88), ack => type_cast_1756_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1622_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1643_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1703_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1734_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1451_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1451_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom52_1745_resized : std_logic_vector(13 downto 0);
    signal R_idxprom52_1745_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1714_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1714_scaled : std_logic_vector(13 downto 0);
    signal add16_1583 : std_logic_vector(31 downto 0);
    signal add27_1598 : std_logic_vector(31 downto 0);
    signal add42_1655 : std_logic_vector(31 downto 0);
    signal add44_1690 : std_logic_vector(31 downto 0);
    signal add57_1763 : std_logic_vector(31 downto 0);
    signal add8_1685 : std_logic_vector(31 downto 0);
    signal add_1568 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1715_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1715_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1715_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1715_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1715_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1715_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1746_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1746_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1746_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1746_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1746_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1746_root_address : std_logic_vector(13 downto 0);
    signal arrayidx53_1748 : std_logic_vector(31 downto 0);
    signal arrayidx_1717 : std_logic_vector(31 downto 0);
    signal call_1398 : std_logic_vector(15 downto 0);
    signal cmp68_1799 : std_logic_vector(0 downto 0);
    signal cmp77_1825 : std_logic_vector(0 downto 0);
    signal cmp_1768 : std_logic_vector(0 downto 0);
    signal conv13_1437 : std_logic_vector(31 downto 0);
    signal conv18_1456 : std_logic_vector(31 downto 0);
    signal conv24_1470 : std_logic_vector(31 downto 0);
    signal conv37_1624 : std_logic_vector(31 downto 0);
    signal conv3_1553 : std_logic_vector(31 downto 0);
    signal conv40_1645 : std_logic_vector(31 downto 0);
    signal conv56_1757 : std_logic_vector(31 downto 0);
    signal conv66_1794 : std_logic_vector(31 downto 0);
    signal conv6_1558 : std_logic_vector(31 downto 0);
    signal conv74_1820 : std_logic_vector(31 downto 0);
    signal conv90_1680 : std_logic_vector(31 downto 0);
    signal div76_1530 : std_logic_vector(31 downto 0);
    signal div_1512 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1520 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1407 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1419 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1429 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1445 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1462 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1478 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1490 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1502 : std_logic_vector(31 downto 0);
    signal idxprom52_1741 : std_logic_vector(63 downto 0);
    signal idxprom_1710 : std_logic_vector(63 downto 0);
    signal inc72_1803 : std_logic_vector(15 downto 0);
    signal inc72x_xinput_dim0x_x2_1808 : std_logic_vector(15 downto 0);
    signal inc_1789 : std_logic_vector(15 downto 0);
    signal indvar_1663 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1781 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1540 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1533 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1815 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1676 : std_logic_vector(15 downto 0);
    signal mul14_1578 : std_logic_vector(31 downto 0);
    signal mul25_1593 : std_logic_vector(31 downto 0);
    signal mul41_1650 : std_logic_vector(31 downto 0);
    signal mul43_1660 : std_logic_vector(31 downto 0);
    signal mul7_1573 : std_logic_vector(31 downto 0);
    signal mul_1563 : std_logic_vector(31 downto 0);
    signal ptr_deref_1410_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1410_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1410_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1410_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1410_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1422_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1422_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1422_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1422_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1422_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1432_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1432_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1432_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1432_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1432_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1448_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1448_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1448_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1448_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1448_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1465_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1465_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1465_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1465_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1465_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1481_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1481_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1481_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1481_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1481_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1493_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1493_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1493_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1493_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1493_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1505_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1505_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1505_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1505_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1505_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1523_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1523_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1523_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1523_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1523_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1720_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1720_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1720_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1720_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1720_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1750_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1750_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1750_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1750_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1750_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1750_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext91_1636 : std_logic_vector(31 downto 0);
    signal sext93_1696 : std_logic_vector(31 downto 0);
    signal sext94_1727 : std_logic_vector(31 downto 0);
    signal sext_1615 : std_logic_vector(31 downto 0);
    signal shr51_1736 : std_logic_vector(31 downto 0);
    signal shr_1705 : std_logic_vector(31 downto 0);
    signal sub19_1630 : std_logic_vector(31 downto 0);
    signal sub30_1603 : std_logic_vector(31 downto 0);
    signal sub31_1609 : std_logic_vector(31 downto 0);
    signal sub_1588 : std_logic_vector(31 downto 0);
    signal tmp12_1433 : std_logic_vector(15 downto 0);
    signal tmp15_1449 : std_logic_vector(31 downto 0);
    signal tmp17_1452 : std_logic_vector(15 downto 0);
    signal tmp1_1411 : std_logic_vector(31 downto 0);
    signal tmp23_1466 : std_logic_vector(15 downto 0);
    signal tmp26_1482 : std_logic_vector(31 downto 0);
    signal tmp35_1494 : std_logic_vector(31 downto 0);
    signal tmp38_1506 : std_logic_vector(31 downto 0);
    signal tmp48_1721 : std_logic_vector(63 downto 0);
    signal tmp4_1423 : std_logic_vector(31 downto 0);
    signal tmp75_1524 : std_logic_vector(31 downto 0);
    signal type_cast_1510_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1528_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1537_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1539_wire : std_logic_vector(15 downto 0);
    signal type_cast_1544_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1546_wire : std_logic_vector(15 downto 0);
    signal type_cast_1551_wire : std_logic_vector(31 downto 0);
    signal type_cast_1556_wire : std_logic_vector(31 downto 0);
    signal type_cast_1607_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1613_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1618_wire : std_logic_vector(31 downto 0);
    signal type_cast_1621_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1628_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1634_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1639_wire : std_logic_vector(31 downto 0);
    signal type_cast_1642_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1667_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1669_wire : std_logic_vector(15 downto 0);
    signal type_cast_1674_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1694_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1699_wire : std_logic_vector(31 downto 0);
    signal type_cast_1702_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1708_wire : std_logic_vector(63 downto 0);
    signal type_cast_1725_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1730_wire : std_logic_vector(31 downto 0);
    signal type_cast_1733_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1739_wire : std_logic_vector(63 downto 0);
    signal type_cast_1755_wire : std_logic_vector(31 downto 0);
    signal type_cast_1761_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1779_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1787_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1792_wire : std_logic_vector(31 downto 0);
    signal type_cast_1812_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1818_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1451_word_address_0 <= "0";
    array_obj_ref_1715_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1715_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1715_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1715_resized_base_address <= "00000000000000";
    array_obj_ref_1746_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1746_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1746_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1746_resized_base_address <= "00000000000000";
    iNsTr_10_1520 <= "00000000000000000000000000000010";
    iNsTr_2_1407 <= "00000000000000000000000000000100";
    iNsTr_3_1419 <= "00000000000000000000000000000011";
    iNsTr_4_1429 <= "00000000000000000000000000000000";
    iNsTr_5_1445 <= "00000000000000000000000000000011";
    iNsTr_6_1462 <= "00000000000000000000000000000001";
    iNsTr_7_1478 <= "00000000000000000000000000000100";
    iNsTr_8_1490 <= "00000000000000000000000000000100";
    iNsTr_9_1502 <= "00000000000000000000000000000011";
    ptr_deref_1410_word_offset_0 <= "0000000";
    ptr_deref_1422_word_offset_0 <= "0000000";
    ptr_deref_1432_word_offset_0 <= "0";
    ptr_deref_1448_word_offset_0 <= "0000000";
    ptr_deref_1465_word_offset_0 <= "0";
    ptr_deref_1481_word_offset_0 <= "0000000";
    ptr_deref_1493_word_offset_0 <= "0000000";
    ptr_deref_1505_word_offset_0 <= "0000000";
    ptr_deref_1523_word_offset_0 <= "0000000";
    ptr_deref_1720_word_offset_0 <= "00000000000000";
    ptr_deref_1750_word_offset_0 <= "00000000000000";
    type_cast_1510_wire_constant <= "00000000000000000000000000000001";
    type_cast_1528_wire_constant <= "00000000000000000000000000000001";
    type_cast_1537_wire_constant <= "0000000000000000";
    type_cast_1544_wire_constant <= "0000000000000000";
    type_cast_1607_wire_constant <= "00000000000000000000000000010000";
    type_cast_1613_wire_constant <= "11111111111111110000000000000000";
    type_cast_1621_wire_constant <= "00000000000000000000000000010000";
    type_cast_1628_wire_constant <= "00000000000000000000000000010000";
    type_cast_1634_wire_constant <= "11111111111111110000000000000000";
    type_cast_1642_wire_constant <= "00000000000000000000000000010000";
    type_cast_1667_wire_constant <= "0000000000000000";
    type_cast_1674_wire_constant <= "0000000000000100";
    type_cast_1694_wire_constant <= "00000000000000000000000000010000";
    type_cast_1702_wire_constant <= "00000000000000000000000000010010";
    type_cast_1725_wire_constant <= "00000000000000000000000000010000";
    type_cast_1733_wire_constant <= "00000000000000000000000000010010";
    type_cast_1761_wire_constant <= "00000000000000000000000000000100";
    type_cast_1779_wire_constant <= "0000000000000001";
    type_cast_1787_wire_constant <= "0000000000000001";
    type_cast_1812_wire_constant <= "0000000000000000";
    phi_stmt_1533: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1537_wire_constant & type_cast_1539_wire;
      req <= phi_stmt_1533_req_0 & phi_stmt_1533_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1533",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1533_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1533,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1533
    phi_stmt_1540: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1544_wire_constant & type_cast_1546_wire;
      req <= phi_stmt_1540_req_0 & phi_stmt_1540_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1540",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1540_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1540,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1540
    phi_stmt_1663: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1667_wire_constant & type_cast_1669_wire;
      req <= phi_stmt_1663_req_0 & phi_stmt_1663_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1663",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1663_ack_0,
          idata => idata,
          odata => indvar_1663,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1663
    -- flow-through select operator MUX_1814_inst
    input_dim1x_x2_1815 <= type_cast_1812_wire_constant when (cmp68_1799(0) /=  '0') else inc_1789;
    addr_of_1716_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1716_final_reg_req_0;
      addr_of_1716_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1716_final_reg_req_1;
      addr_of_1716_final_reg_ack_1<= rack(0);
      addr_of_1716_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1716_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1715_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1717,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1747_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1747_final_reg_req_0;
      addr_of_1747_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1747_final_reg_req_1;
      addr_of_1747_final_reg_ack_1<= rack(0);
      addr_of_1747_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1747_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1746_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx53_1748,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1436_inst_req_0;
      type_cast_1436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1436_inst_req_1;
      type_cast_1436_inst_ack_1<= rack(0);
      type_cast_1436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_1433,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_1437,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1455_inst_req_0;
      type_cast_1455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1455_inst_req_1;
      type_cast_1455_inst_ack_1<= rack(0);
      type_cast_1455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp17_1452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_1456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1469_inst_req_0;
      type_cast_1469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1469_inst_req_1;
      type_cast_1469_inst_ack_1<= rack(0);
      type_cast_1469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp23_1466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_1470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1539_inst_req_0;
      type_cast_1539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1539_inst_req_1;
      type_cast_1539_inst_ack_1<= rack(0);
      type_cast_1539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1539_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1546_inst_req_0;
      type_cast_1546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1546_inst_req_1;
      type_cast_1546_inst_ack_1<= rack(0);
      type_cast_1546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1546_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc72x_xinput_dim0x_x2_1808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1546_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1552_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1552_inst_req_0;
      type_cast_1552_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1552_inst_req_1;
      type_cast_1552_inst_ack_1<= rack(0);
      type_cast_1552_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1552_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1551_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1553,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1557_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1557_inst_req_0;
      type_cast_1557_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1557_inst_req_1;
      type_cast_1557_inst_ack_1<= rack(0);
      type_cast_1557_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1557_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1556_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv6_1558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1618_inst
    process(sext_1615) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1615(31 downto 0);
      type_cast_1618_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1623_inst
    process(ASHR_i32_i32_1622_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1622_wire(31 downto 0);
      conv37_1624 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1639_inst
    process(sext91_1636) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext91_1636(31 downto 0);
      type_cast_1639_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1644_inst
    process(ASHR_i32_i32_1643_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1643_wire(31 downto 0);
      conv40_1645 <= tmp_var; -- 
    end process;
    type_cast_1669_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1669_inst_req_0;
      type_cast_1669_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1669_inst_req_1;
      type_cast_1669_inst_ack_1<= rack(0);
      type_cast_1669_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1669_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1669_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1679_inst_req_0;
      type_cast_1679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1679_inst_req_1;
      type_cast_1679_inst_ack_1<= rack(0);
      type_cast_1679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1680,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1699_inst
    process(sext93_1696) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext93_1696(31 downto 0);
      type_cast_1699_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1704_inst
    process(ASHR_i32_i32_1703_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1703_wire(31 downto 0);
      shr_1705 <= tmp_var; -- 
    end process;
    type_cast_1709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1709_inst_req_0;
      type_cast_1709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1709_inst_req_1;
      type_cast_1709_inst_ack_1<= rack(0);
      type_cast_1709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1708_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1730_inst
    process(sext94_1727) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext94_1727(31 downto 0);
      type_cast_1730_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1735_inst
    process(ASHR_i32_i32_1734_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1734_wire(31 downto 0);
      shr51_1736 <= tmp_var; -- 
    end process;
    type_cast_1740_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1740_inst_req_0;
      type_cast_1740_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1740_inst_req_1;
      type_cast_1740_inst_ack_1<= rack(0);
      type_cast_1740_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1740_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1739_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom52_1741,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1756_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1756_inst_req_0;
      type_cast_1756_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1756_inst_req_1;
      type_cast_1756_inst_ack_1<= rack(0);
      type_cast_1756_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1756_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1755_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1793_inst_req_0;
      type_cast_1793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1793_inst_req_1;
      type_cast_1793_inst_ack_1<= rack(0);
      type_cast_1793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1792_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1802_inst_req_0;
      type_cast_1802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1802_inst_req_1;
      type_cast_1802_inst_ack_1<= rack(0);
      type_cast_1802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp68_1799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc72_1803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1819_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1819_inst_req_0;
      type_cast_1819_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1819_inst_req_1;
      type_cast_1819_inst_ack_1<= rack(0);
      type_cast_1819_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1819_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1818_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_1820,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1451_gather_scatter
    process(LOAD_padding_1451_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1451_data_0;
      ov(15 downto 0) := iv;
      tmp17_1452 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1715_index_1_rename
    process(R_idxprom_1714_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1714_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1714_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1715_index_1_resize
    process(idxprom_1710) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1710;
      ov := iv(13 downto 0);
      R_idxprom_1714_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1715_root_address_inst
    process(array_obj_ref_1715_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1715_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1715_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1746_index_1_rename
    process(R_idxprom52_1745_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom52_1745_resized;
      ov(13 downto 0) := iv;
      R_idxprom52_1745_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1746_index_1_resize
    process(idxprom52_1741) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom52_1741;
      ov := iv(13 downto 0);
      R_idxprom52_1745_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1746_root_address_inst
    process(array_obj_ref_1746_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1746_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1746_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1410_addr_0
    process(ptr_deref_1410_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1410_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1410_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1410_base_resize
    process(iNsTr_2_1407) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1407;
      ov := iv(6 downto 0);
      ptr_deref_1410_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1410_gather_scatter
    process(ptr_deref_1410_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1410_data_0;
      ov(31 downto 0) := iv;
      tmp1_1411 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1410_root_address_inst
    process(ptr_deref_1410_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1410_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1410_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1422_addr_0
    process(ptr_deref_1422_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1422_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1422_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1422_base_resize
    process(iNsTr_3_1419) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1419;
      ov := iv(6 downto 0);
      ptr_deref_1422_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1422_gather_scatter
    process(ptr_deref_1422_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1422_data_0;
      ov(31 downto 0) := iv;
      tmp4_1423 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1422_root_address_inst
    process(ptr_deref_1422_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1422_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1422_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1432_addr_0
    process(ptr_deref_1432_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1432_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1432_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1432_base_resize
    process(iNsTr_4_1429) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1429;
      ov := iv(0 downto 0);
      ptr_deref_1432_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1432_gather_scatter
    process(ptr_deref_1432_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1432_data_0;
      ov(15 downto 0) := iv;
      tmp12_1433 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1432_root_address_inst
    process(ptr_deref_1432_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1432_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1432_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1448_addr_0
    process(ptr_deref_1448_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1448_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1448_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1448_base_resize
    process(iNsTr_5_1445) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1445;
      ov := iv(6 downto 0);
      ptr_deref_1448_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1448_gather_scatter
    process(ptr_deref_1448_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1448_data_0;
      ov(31 downto 0) := iv;
      tmp15_1449 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1448_root_address_inst
    process(ptr_deref_1448_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1448_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1448_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1465_addr_0
    process(ptr_deref_1465_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1465_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1465_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1465_base_resize
    process(iNsTr_6_1462) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1462;
      ov := iv(0 downto 0);
      ptr_deref_1465_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1465_gather_scatter
    process(ptr_deref_1465_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1465_data_0;
      ov(15 downto 0) := iv;
      tmp23_1466 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1465_root_address_inst
    process(ptr_deref_1465_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1465_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1465_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1481_addr_0
    process(ptr_deref_1481_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1481_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1481_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1481_base_resize
    process(iNsTr_7_1478) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1478;
      ov := iv(6 downto 0);
      ptr_deref_1481_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1481_gather_scatter
    process(ptr_deref_1481_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1481_data_0;
      ov(31 downto 0) := iv;
      tmp26_1482 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1481_root_address_inst
    process(ptr_deref_1481_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1481_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1481_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1493_addr_0
    process(ptr_deref_1493_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1493_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1493_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1493_base_resize
    process(iNsTr_8_1490) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1490;
      ov := iv(6 downto 0);
      ptr_deref_1493_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1493_gather_scatter
    process(ptr_deref_1493_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1493_data_0;
      ov(31 downto 0) := iv;
      tmp35_1494 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1493_root_address_inst
    process(ptr_deref_1493_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1493_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1493_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1505_addr_0
    process(ptr_deref_1505_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1505_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1505_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1505_base_resize
    process(iNsTr_9_1502) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1502;
      ov := iv(6 downto 0);
      ptr_deref_1505_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1505_gather_scatter
    process(ptr_deref_1505_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1505_data_0;
      ov(31 downto 0) := iv;
      tmp38_1506 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1505_root_address_inst
    process(ptr_deref_1505_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1505_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1505_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1523_addr_0
    process(ptr_deref_1523_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1523_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1523_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1523_base_resize
    process(iNsTr_10_1520) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1520;
      ov := iv(6 downto 0);
      ptr_deref_1523_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1523_gather_scatter
    process(ptr_deref_1523_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1523_data_0;
      ov(31 downto 0) := iv;
      tmp75_1524 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1523_root_address_inst
    process(ptr_deref_1523_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1523_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1523_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_addr_0
    process(ptr_deref_1720_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1720_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1720_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_base_resize
    process(arrayidx_1717) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1717;
      ov := iv(13 downto 0);
      ptr_deref_1720_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_gather_scatter
    process(ptr_deref_1720_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1720_data_0;
      ov(63 downto 0) := iv;
      tmp48_1721 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_root_address_inst
    process(ptr_deref_1720_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1720_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1720_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1750_addr_0
    process(ptr_deref_1750_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1750_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1750_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1750_base_resize
    process(arrayidx53_1748) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx53_1748;
      ov := iv(13 downto 0);
      ptr_deref_1750_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1750_gather_scatter
    process(tmp48_1721) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp48_1721;
      ov(63 downto 0) := iv;
      ptr_deref_1750_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1750_root_address_inst
    process(ptr_deref_1750_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1750_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1750_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1769_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1768;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1769_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1769_branch_req_0,
          ack0 => if_stmt_1769_branch_ack_0,
          ack1 => if_stmt_1769_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1826_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1825;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1826_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1826_branch_req_0,
          ack0 => if_stmt_1826_branch_ack_0,
          ack1 => if_stmt_1826_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1780_inst
    process(indvar_1663) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1663, type_cast_1779_wire_constant, tmp_var);
      indvarx_xnext_1781 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1788_inst
    process(input_dim1x_x1x_xph_1533) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1533, type_cast_1787_wire_constant, tmp_var);
      inc_1789 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1807_inst
    process(inc72_1803, input_dim0x_x2x_xph_1540) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc72_1803, input_dim0x_x2x_xph_1540, tmp_var);
      inc72x_xinput_dim0x_x2_1808 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1567_inst
    process(mul_1563, conv3_1553) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1563, conv3_1553, tmp_var);
      add_1568 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1582_inst
    process(mul14_1578, tmp15_1449) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul14_1578, tmp15_1449, tmp_var);
      add16_1583 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1597_inst
    process(mul25_1593, tmp26_1482) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul25_1593, tmp26_1482, tmp_var);
      add27_1598 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1614_inst
    process(sub31_1609) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub31_1609, type_cast_1613_wire_constant, tmp_var);
      sext_1615 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1635_inst
    process(sub19_1630) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub19_1630, type_cast_1634_wire_constant, tmp_var);
      sext91_1636 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1654_inst
    process(conv37_1624, mul41_1650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv37_1624, mul41_1650, tmp_var);
      add42_1655 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1684_inst
    process(mul7_1573, conv90_1680) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul7_1573, conv90_1680, tmp_var);
      add8_1685 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1689_inst
    process(mul43_1660, conv90_1680) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul43_1660, conv90_1680, tmp_var);
      add44_1690 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1762_inst
    process(conv56_1757) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv56_1757, type_cast_1761_wire_constant, tmp_var);
      add57_1763 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1622_inst
    process(type_cast_1618_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1618_wire, type_cast_1621_wire_constant, tmp_var);
      ASHR_i32_i32_1622_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1643_inst
    process(type_cast_1639_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1639_wire, type_cast_1642_wire_constant, tmp_var);
      ASHR_i32_i32_1643_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1703_inst
    process(type_cast_1699_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1699_wire, type_cast_1702_wire_constant, tmp_var);
      ASHR_i32_i32_1703_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1734_inst
    process(type_cast_1730_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1730_wire, type_cast_1733_wire_constant, tmp_var);
      ASHR_i32_i32_1734_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1798_inst
    process(conv66_1794, div_1512) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv66_1794, div_1512, tmp_var);
      cmp68_1799 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1824_inst
    process(conv74_1820, div76_1530) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv74_1820, div76_1530, tmp_var);
      cmp77_1825 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1511_inst
    process(tmp4_1423) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1423, type_cast_1510_wire_constant, tmp_var);
      div_1512 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1529_inst
    process(tmp75_1524) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp75_1524, type_cast_1528_wire_constant, tmp_var);
      div76_1530 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1675_inst
    process(indvar_1663) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1663, type_cast_1674_wire_constant, tmp_var);
      input_dim2x_x1_1676 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1562_inst
    process(tmp4_1423, conv6_1558) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp4_1423, conv6_1558, tmp_var);
      mul_1563 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1572_inst
    process(add_1568, tmp1_1411) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1568, tmp1_1411, tmp_var);
      mul7_1573 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1577_inst
    process(conv13_1437, conv6_1558) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv13_1437, conv6_1558, tmp_var);
      mul14_1578 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1592_inst
    process(conv24_1470, conv3_1553) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv24_1470, conv3_1553, tmp_var);
      mul25_1593 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1649_inst
    process(tmp38_1506, conv40_1645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp38_1506, conv40_1645, tmp_var);
      mul41_1650 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1659_inst
    process(add42_1655, tmp35_1494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add42_1655, tmp35_1494, tmp_var);
      mul43_1660 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1608_inst
    process(sub30_1603) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub30_1603, type_cast_1607_wire_constant, tmp_var);
      sub31_1609 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1629_inst
    process(sub_1588) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_1588, type_cast_1628_wire_constant, tmp_var);
      sub19_1630 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1695_inst
    process(add8_1685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add8_1685, type_cast_1694_wire_constant, tmp_var);
      sext93_1696 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1726_inst
    process(add44_1690) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add44_1690, type_cast_1725_wire_constant, tmp_var);
      sext94_1727 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1587_inst
    process(add16_1583, conv18_1456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add16_1583, conv18_1456, tmp_var);
      sub_1588 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1602_inst
    process(add27_1598, conv18_1456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add27_1598, conv18_1456, tmp_var);
      sub30_1603 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1767_inst
    process(add57_1763, tmp1_1411) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add57_1763, tmp1_1411, tmp_var);
      cmp_1768 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_1715_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1714_scaled;
      array_obj_ref_1715_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1715_index_offset_req_0;
      array_obj_ref_1715_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1715_index_offset_req_1;
      array_obj_ref_1715_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_1746_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom52_1745_scaled;
      array_obj_ref_1746_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1746_index_offset_req_0;
      array_obj_ref_1746_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1746_index_offset_req_1;
      array_obj_ref_1746_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_1551_inst
    process(input_dim1x_x1x_xph_1533) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1533, tmp_var);
      type_cast_1551_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1556_inst
    process(input_dim0x_x2x_xph_1540) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1540, tmp_var);
      type_cast_1556_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1708_inst
    process(shr_1705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1705, tmp_var);
      type_cast_1708_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1739_inst
    process(shr51_1736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr51_1736, tmp_var);
      type_cast_1739_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1755_inst
    process(input_dim2x_x1_1676) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1676, tmp_var);
      type_cast_1755_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1792_inst
    process(inc_1789) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1789, tmp_var);
      type_cast_1792_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1818_inst
    process(inc72x_xinput_dim0x_x2_1808) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc72x_xinput_dim0x_x2_1808, tmp_var);
      type_cast_1818_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1451_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1451_load_0_req_0;
      LOAD_padding_1451_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1451_load_0_req_1;
      LOAD_padding_1451_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1451_word_address_0;
      LOAD_padding_1451_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1523_load_0 ptr_deref_1422_load_0 ptr_deref_1410_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1523_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1422_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1410_load_0_req_0;
      ptr_deref_1523_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1422_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1410_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1523_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1422_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1410_load_0_req_1;
      ptr_deref_1523_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1422_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1410_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1523_word_address_0 & ptr_deref_1422_word_address_0 & ptr_deref_1410_word_address_0;
      ptr_deref_1523_data_0 <= data_out(95 downto 64);
      ptr_deref_1422_data_0 <= data_out(63 downto 32);
      ptr_deref_1410_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1465_load_0 ptr_deref_1432_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1465_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1432_load_0_req_0;
      ptr_deref_1465_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1432_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1465_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1432_load_0_req_1;
      ptr_deref_1465_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1432_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1465_word_address_0 & ptr_deref_1432_word_address_0;
      ptr_deref_1465_data_0 <= data_out(31 downto 16);
      ptr_deref_1432_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1481_load_0 ptr_deref_1448_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1481_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1448_load_0_req_0;
      ptr_deref_1481_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1448_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1481_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1448_load_0_req_1;
      ptr_deref_1481_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1448_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1481_word_address_0 & ptr_deref_1448_word_address_0;
      ptr_deref_1481_data_0 <= data_out(63 downto 32);
      ptr_deref_1448_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1493_load_0 ptr_deref_1505_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1493_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1505_load_0_req_0;
      ptr_deref_1493_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1505_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1493_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1505_load_0_req_1;
      ptr_deref_1493_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1505_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1493_word_address_0 & ptr_deref_1505_word_address_0;
      ptr_deref_1493_data_0 <= data_out(63 downto 32);
      ptr_deref_1505_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1720_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1720_load_0_req_0;
      ptr_deref_1720_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1720_load_0_req_1;
      ptr_deref_1720_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1720_word_address_0;
      ptr_deref_1720_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1750_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1750_store_0_req_0;
      ptr_deref_1750_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1750_store_0_req_1;
      ptr_deref_1750_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1750_word_address_0;
      data_in <= ptr_deref_1750_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1397_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_start_1397_inst_req_0;
      RPIPE_Block0_start_1397_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_start_1397_inst_req_1;
      RPIPE_Block0_start_1397_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1398 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1834_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1834_inst_req_0;
      WPIPE_Block0_done_1834_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1834_inst_req_1;
      WPIPE_Block0_done_1834_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1398;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_5316_start: Boolean;
  signal convTransposeB_CP_5316_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1889_load_0_req_1 : boolean;
  signal ptr_deref_1889_load_0_ack_1 : boolean;
  signal ptr_deref_1879_load_0_req_0 : boolean;
  signal type_cast_1867_inst_req_1 : boolean;
  signal ptr_deref_1889_load_0_ack_0 : boolean;
  signal ptr_deref_1879_load_0_ack_0 : boolean;
  signal ptr_deref_1905_load_0_req_0 : boolean;
  signal type_cast_1867_inst_ack_1 : boolean;
  signal ptr_deref_1905_load_0_ack_0 : boolean;
  signal type_cast_1867_inst_req_0 : boolean;
  signal type_cast_1893_inst_ack_1 : boolean;
  signal type_cast_1893_inst_req_0 : boolean;
  signal type_cast_1867_inst_ack_0 : boolean;
  signal type_cast_1893_inst_ack_0 : boolean;
  signal ptr_deref_1905_load_0_req_1 : boolean;
  signal type_cast_1893_inst_req_1 : boolean;
  signal ptr_deref_1889_load_0_req_0 : boolean;
  signal LOAD_padding_1908_load_0_ack_1 : boolean;
  signal LOAD_padding_1908_load_0_req_1 : boolean;
  signal LOAD_padding_1908_load_0_req_0 : boolean;
  signal LOAD_padding_1908_load_0_ack_0 : boolean;
  signal WPIPE_Block1_done_2305_inst_ack_1 : boolean;
  signal WPIPE_Block1_done_2305_inst_req_1 : boolean;
  signal type_cast_2283_inst_ack_1 : boolean;
  signal ptr_deref_1857_load_0_ack_1 : boolean;
  signal type_cast_1989_inst_ack_0 : boolean;
  signal ptr_deref_1879_load_0_ack_1 : boolean;
  signal ptr_deref_1879_load_0_req_1 : boolean;
  signal ptr_deref_1905_load_0_ack_1 : boolean;
  signal phi_stmt_2280_req_0 : boolean;
  signal if_stmt_2297_branch_ack_1 : boolean;
  signal type_cast_1987_inst_req_1 : boolean;
  signal type_cast_1987_inst_ack_1 : boolean;
  signal phi_stmt_2274_ack_0 : boolean;
  signal phi_stmt_2280_ack_0 : boolean;
  signal phi_stmt_1984_req_0 : boolean;
  signal type_cast_1989_inst_req_1 : boolean;
  signal type_cast_1989_inst_ack_1 : boolean;
  signal type_cast_2279_inst_ack_0 : boolean;
  signal type_cast_2279_inst_req_0 : boolean;
  signal type_cast_2279_inst_req_1 : boolean;
  signal type_cast_2279_inst_ack_1 : boolean;
  signal phi_stmt_2274_req_1 : boolean;
  signal type_cast_2115_inst_req_1 : boolean;
  signal type_cast_2115_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1844_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1844_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1844_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1844_inst_ack_1 : boolean;
  signal ptr_deref_1857_load_0_req_0 : boolean;
  signal ptr_deref_1857_load_0_ack_0 : boolean;
  signal ptr_deref_1857_load_0_req_1 : boolean;
  signal type_cast_1912_inst_req_0 : boolean;
  signal type_cast_1912_inst_ack_0 : boolean;
  signal type_cast_1912_inst_req_1 : boolean;
  signal type_cast_1912_inst_ack_1 : boolean;
  signal ptr_deref_1922_load_0_req_0 : boolean;
  signal ptr_deref_1922_load_0_ack_0 : boolean;
  signal ptr_deref_1922_load_0_req_1 : boolean;
  signal ptr_deref_1922_load_0_ack_1 : boolean;
  signal type_cast_1926_inst_req_0 : boolean;
  signal type_cast_1926_inst_ack_0 : boolean;
  signal type_cast_1926_inst_req_1 : boolean;
  signal type_cast_1926_inst_ack_1 : boolean;
  signal ptr_deref_1938_load_0_req_0 : boolean;
  signal ptr_deref_1938_load_0_ack_0 : boolean;
  signal ptr_deref_1938_load_0_req_1 : boolean;
  signal ptr_deref_1938_load_0_ack_1 : boolean;
  signal ptr_deref_1950_load_0_req_0 : boolean;
  signal ptr_deref_1950_load_0_ack_0 : boolean;
  signal ptr_deref_1950_load_0_req_1 : boolean;
  signal ptr_deref_1950_load_0_ack_1 : boolean;
  signal ptr_deref_1962_load_0_req_0 : boolean;
  signal ptr_deref_1962_load_0_ack_0 : boolean;
  signal ptr_deref_1962_load_0_req_1 : boolean;
  signal ptr_deref_1962_load_0_ack_1 : boolean;
  signal ptr_deref_1974_load_0_req_0 : boolean;
  signal ptr_deref_1974_load_0_ack_0 : boolean;
  signal ptr_deref_1974_load_0_req_1 : boolean;
  signal ptr_deref_1974_load_0_ack_1 : boolean;
  signal type_cast_2001_inst_req_0 : boolean;
  signal type_cast_2001_inst_ack_0 : boolean;
  signal type_cast_2001_inst_req_1 : boolean;
  signal type_cast_2001_inst_ack_1 : boolean;
  signal type_cast_2006_inst_req_0 : boolean;
  signal type_cast_2006_inst_ack_0 : boolean;
  signal type_cast_2006_inst_req_1 : boolean;
  signal type_cast_2006_inst_ack_1 : boolean;
  signal WPIPE_Block1_done_2305_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2305_inst_req_0 : boolean;
  signal type_cast_1989_inst_req_0 : boolean;
  signal type_cast_2128_inst_req_0 : boolean;
  signal type_cast_2128_inst_ack_0 : boolean;
  signal type_cast_2128_inst_req_1 : boolean;
  signal type_cast_2128_inst_ack_1 : boolean;
  signal type_cast_2283_inst_req_1 : boolean;
  signal type_cast_2158_inst_req_0 : boolean;
  signal type_cast_2158_inst_ack_0 : boolean;
  signal type_cast_2115_inst_ack_0 : boolean;
  signal type_cast_2158_inst_req_1 : boolean;
  signal type_cast_2158_inst_ack_1 : boolean;
  signal phi_stmt_2274_req_0 : boolean;
  signal type_cast_2277_inst_ack_1 : boolean;
  signal type_cast_2277_inst_req_1 : boolean;
  signal type_cast_2277_inst_ack_0 : boolean;
  signal type_cast_2115_inst_req_0 : boolean;
  signal array_obj_ref_2164_index_offset_req_0 : boolean;
  signal array_obj_ref_2164_index_offset_ack_0 : boolean;
  signal array_obj_ref_2164_index_offset_req_1 : boolean;
  signal array_obj_ref_2164_index_offset_ack_1 : boolean;
  signal phi_stmt_1990_req_0 : boolean;
  signal addr_of_2165_final_reg_req_0 : boolean;
  signal addr_of_2165_final_reg_ack_0 : boolean;
  signal addr_of_2165_final_reg_req_1 : boolean;
  signal addr_of_2165_final_reg_ack_1 : boolean;
  signal type_cast_2277_inst_req_0 : boolean;
  signal phi_stmt_1990_req_1 : boolean;
  signal type_cast_1987_inst_ack_0 : boolean;
  signal ptr_deref_2169_load_0_req_0 : boolean;
  signal ptr_deref_2169_load_0_ack_0 : boolean;
  signal ptr_deref_2169_load_0_req_1 : boolean;
  signal ptr_deref_2169_load_0_ack_1 : boolean;
  signal type_cast_1996_inst_ack_1 : boolean;
  signal if_stmt_2297_branch_req_0 : boolean;
  signal type_cast_1996_inst_req_1 : boolean;
  signal type_cast_2189_inst_req_0 : boolean;
  signal type_cast_2189_inst_ack_0 : boolean;
  signal type_cast_2189_inst_req_1 : boolean;
  signal type_cast_2189_inst_ack_1 : boolean;
  signal phi_stmt_2280_req_1 : boolean;
  signal type_cast_2285_inst_ack_1 : boolean;
  signal type_cast_1996_inst_ack_0 : boolean;
  signal type_cast_1996_inst_req_0 : boolean;
  signal array_obj_ref_2195_index_offset_req_0 : boolean;
  signal array_obj_ref_2195_index_offset_ack_0 : boolean;
  signal array_obj_ref_2195_index_offset_req_1 : boolean;
  signal array_obj_ref_2195_index_offset_ack_1 : boolean;
  signal phi_stmt_2112_ack_0 : boolean;
  signal addr_of_2196_final_reg_req_0 : boolean;
  signal addr_of_2196_final_reg_ack_0 : boolean;
  signal addr_of_2196_final_reg_req_1 : boolean;
  signal phi_stmt_2112_req_1 : boolean;
  signal addr_of_2196_final_reg_ack_1 : boolean;
  signal type_cast_2285_inst_req_1 : boolean;
  signal type_cast_2285_inst_ack_0 : boolean;
  signal type_cast_2285_inst_req_0 : boolean;
  signal type_cast_1987_inst_req_0 : boolean;
  signal ptr_deref_2199_store_0_req_0 : boolean;
  signal ptr_deref_2199_store_0_ack_0 : boolean;
  signal ptr_deref_2199_store_0_req_1 : boolean;
  signal ptr_deref_2199_store_0_ack_1 : boolean;
  signal type_cast_2205_inst_req_0 : boolean;
  signal type_cast_2205_inst_ack_0 : boolean;
  signal type_cast_2205_inst_req_1 : boolean;
  signal type_cast_2205_inst_ack_1 : boolean;
  signal if_stmt_2218_branch_req_0 : boolean;
  signal if_stmt_2218_branch_ack_1 : boolean;
  signal if_stmt_2218_branch_ack_0 : boolean;
  signal type_cast_2283_inst_ack_0 : boolean;
  signal if_stmt_2297_branch_ack_0 : boolean;
  signal phi_stmt_1990_ack_0 : boolean;
  signal phi_stmt_1984_ack_0 : boolean;
  signal type_cast_2242_inst_req_0 : boolean;
  signal type_cast_2242_inst_ack_0 : boolean;
  signal type_cast_2242_inst_req_1 : boolean;
  signal phi_stmt_2112_req_0 : boolean;
  signal type_cast_2242_inst_ack_1 : boolean;
  signal type_cast_2283_inst_req_0 : boolean;
  signal if_stmt_2249_branch_req_0 : boolean;
  signal phi_stmt_1984_req_1 : boolean;
  signal if_stmt_2249_branch_ack_1 : boolean;
  signal if_stmt_2249_branch_ack_0 : boolean;
  signal type_cast_2270_inst_req_0 : boolean;
  signal type_cast_2270_inst_ack_0 : boolean;
  signal type_cast_2270_inst_req_1 : boolean;
  signal type_cast_2270_inst_ack_1 : boolean;
  signal type_cast_2290_inst_req_0 : boolean;
  signal type_cast_2290_inst_ack_0 : boolean;
  signal type_cast_2290_inst_req_1 : boolean;
  signal type_cast_2290_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_5316_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5316_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_5316_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5316_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_5316: Block -- control-path 
    signal convTransposeB_CP_5316_elements: BooleanArray(112 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_5316_elements(0) <= convTransposeB_CP_5316_start;
    convTransposeB_CP_5316_symbol <= convTransposeB_CP_5316_elements(72);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1842/$entry
      -- CP-element group 0: 	 branch_block_stmt_1842/branch_block_stmt_1842__entry__
      -- CP-element group 0: 	 branch_block_stmt_1842/assign_stmt_1845__entry__
      -- CP-element group 0: 	 branch_block_stmt_1842/assign_stmt_1845/$entry
      -- CP-element group 0: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_Sample/rr
      -- 
    rr_5374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(0), ack => RPIPE_Block1_start_1844_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_Update/cr
      -- 
    ra_5375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1844_inst_ack_0, ack => convTransposeB_CP_5316_elements(1)); -- 
    cr_5379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(1), ack => RPIPE_Block1_start_1844_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1845__exit__
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981__entry__
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1845/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1845/RPIPE_Block1_start_1844_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/word_access_complete/word_0/cr
      -- 
    ca_5380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1844_inst_ack_1, ack => convTransposeB_CP_5316_elements(2)); -- 
    cr_5541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1889_load_0_req_1); -- 
    rr_5480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1879_load_0_req_0); -- 
    cr_5446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => type_cast_1867_inst_req_1); -- 
    rr_5594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1905_load_0_req_0); -- 
    cr_5605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1905_load_0_req_1); -- 
    cr_5560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => type_cast_1893_inst_req_1); -- 
    rr_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1889_load_0_req_0); -- 
    cr_5638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => LOAD_padding_1908_load_0_req_1); -- 
    rr_5627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => LOAD_padding_1908_load_0_req_0); -- 
    cr_5491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1879_load_0_req_1); -- 
    rr_5416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1857_load_0_req_0); -- 
    cr_5427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1857_load_0_req_1); -- 
    cr_5657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => type_cast_1912_inst_req_1); -- 
    rr_5691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1922_load_0_req_0); -- 
    cr_5702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1922_load_0_req_1); -- 
    cr_5721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => type_cast_1926_inst_req_1); -- 
    rr_5755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1938_load_0_req_0); -- 
    cr_5766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1938_load_0_req_1); -- 
    rr_5805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1950_load_0_req_0); -- 
    cr_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1950_load_0_req_1); -- 
    rr_5855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1962_load_0_req_0); -- 
    cr_5866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1962_load_0_req_1); -- 
    rr_5905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1974_load_0_req_0); -- 
    cr_5916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(2), ack => ptr_deref_1974_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Sample/word_access_start/word_0/ra
      -- 
    ra_5417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1857_load_0_ack_0, ack => convTransposeB_CP_5316_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/ptr_deref_1857_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/ptr_deref_1857_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/ptr_deref_1857_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/ptr_deref_1857_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1857_Update/word_access_complete/word_0/$exit
      -- 
    ca_5428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1857_load_0_ack_1, ack => convTransposeB_CP_5316_elements(4)); -- 
    rr_5441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(4), ack => type_cast_1867_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_sample_completed_
      -- 
    ra_5442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_0, ack => convTransposeB_CP_5316_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1867_Update/ca
      -- 
    ca_5447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_1, ack => convTransposeB_CP_5316_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Sample/$exit
      -- 
    ra_5481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1879_load_0_ack_0, ack => convTransposeB_CP_5316_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/ptr_deref_1879_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/ptr_deref_1879_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/ptr_deref_1879_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/ptr_deref_1879_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1879_Update/word_access_complete/word_0/ca
      -- 
    ca_5492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1879_load_0_ack_1, ack => convTransposeB_CP_5316_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Sample/$exit
      -- 
    ra_5531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1889_load_0_ack_0, ack => convTransposeB_CP_5316_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/ptr_deref_1889_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/ptr_deref_1889_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/ptr_deref_1889_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1889_Update/ptr_deref_1889_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_sample_start_
      -- 
    ca_5542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1889_load_0_ack_1, ack => convTransposeB_CP_5316_elements(10)); -- 
    rr_5555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(10), ack => type_cast_1893_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_sample_completed_
      -- 
    ra_5556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1893_inst_ack_0, ack => convTransposeB_CP_5316_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1893_update_completed_
      -- 
    ca_5561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1893_inst_ack_1, ack => convTransposeB_CP_5316_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Sample/word_access_start/$exit
      -- 
    ra_5595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_0, ack => convTransposeB_CP_5316_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/ptr_deref_1905_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/ptr_deref_1905_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/ptr_deref_1905_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1905_Update/ptr_deref_1905_Merge/$entry
      -- 
    ca_5606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_1, ack => convTransposeB_CP_5316_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_sample_completed_
      -- 
    ra_5628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1908_load_0_ack_0, ack => convTransposeB_CP_5316_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (12) 
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/LOAD_padding_1908_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/LOAD_padding_1908_Merge/merge_ack
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/LOAD_padding_1908_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/LOAD_padding_1908_Update/LOAD_padding_1908_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_Sample/rr
      -- 
    ca_5639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1908_load_0_ack_1, ack => convTransposeB_CP_5316_elements(16)); -- 
    rr_5652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(16), ack => type_cast_1912_inst_req_0); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_Sample/ra
      -- 
    ra_5653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1912_inst_ack_0, ack => convTransposeB_CP_5316_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	31 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1912_Update/ca
      -- 
    ca_5658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1912_inst_ack_1, ack => convTransposeB_CP_5316_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Sample/word_access_start/word_0/ra
      -- 
    ra_5692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1922_load_0_ack_0, ack => convTransposeB_CP_5316_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/ptr_deref_1922_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/ptr_deref_1922_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/ptr_deref_1922_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1922_Update/ptr_deref_1922_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_Sample/rr
      -- 
    ca_5703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1922_load_0_ack_1, ack => convTransposeB_CP_5316_elements(20)); -- 
    rr_5716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(20), ack => type_cast_1926_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_Sample/ra
      -- 
    ra_5717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1926_inst_ack_0, ack => convTransposeB_CP_5316_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/type_cast_1926_Update/ca
      -- 
    ca_5722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1926_inst_ack_1, ack => convTransposeB_CP_5316_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Sample/word_access_start/word_0/ra
      -- 
    ra_5756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1938_load_0_ack_0, ack => convTransposeB_CP_5316_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/ptr_deref_1938_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/ptr_deref_1938_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/ptr_deref_1938_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1938_Update/ptr_deref_1938_Merge/merge_ack
      -- 
    ca_5767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1938_load_0_ack_1, ack => convTransposeB_CP_5316_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Sample/word_access_start/word_0/ra
      -- 
    ra_5806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1950_load_0_ack_0, ack => convTransposeB_CP_5316_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/ptr_deref_1950_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/ptr_deref_1950_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/ptr_deref_1950_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1950_Update/ptr_deref_1950_Merge/merge_ack
      -- 
    ca_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1950_load_0_ack_1, ack => convTransposeB_CP_5316_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Sample/word_access_start/word_0/ra
      -- 
    ra_5856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1962_load_0_ack_0, ack => convTransposeB_CP_5316_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/ptr_deref_1962_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/ptr_deref_1962_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/ptr_deref_1962_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1962_Update/ptr_deref_1962_Merge/merge_ack
      -- 
    ca_5867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1962_load_0_ack_1, ack => convTransposeB_CP_5316_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Sample/word_access_start/word_0/ra
      -- 
    ra_5906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1974_load_0_ack_0, ack => convTransposeB_CP_5316_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/ptr_deref_1974_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/ptr_deref_1974_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/ptr_deref_1974_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/ptr_deref_1974_Update/ptr_deref_1974_Merge/merge_ack
      -- 
    ca_5917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1974_load_0_ack_1, ack => convTransposeB_CP_5316_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	18 
    -- CP-element group 31: 	6 
    -- CP-element group 31: 	8 
    -- CP-element group 31: 	12 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	73 
    -- CP-element group 31: 	74 
    -- CP-element group 31: 	75 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/$entry
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/$entry
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981__exit__
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1842/assign_stmt_1854_to_assign_stmt_1981/$exit
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/$entry
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Sample/$entry
      -- 
    cr_6364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(31), ack => type_cast_1987_inst_req_1); -- 
    rr_6359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(31), ack => type_cast_1987_inst_req_0); -- 
    convTransposeB_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(22) & convTransposeB_CP_5316_elements(24) & convTransposeB_CP_5316_elements(14) & convTransposeB_CP_5316_elements(26) & convTransposeB_CP_5316_elements(28) & convTransposeB_CP_5316_elements(30) & convTransposeB_CP_5316_elements(18) & convTransposeB_CP_5316_elements(6) & convTransposeB_CP_5316_elements(8) & convTransposeB_CP_5316_elements(12);
      gj_convTransposeB_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	88 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_Sample/ra
      -- 
    ra_5934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2001_inst_ack_0, ack => convTransposeB_CP_5316_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	88 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_Update/ca
      -- 
    ca_5939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2001_inst_ack_1, ack => convTransposeB_CP_5316_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	88 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_Sample/ra
      -- 
    ra_5948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2006_inst_ack_0, ack => convTransposeB_CP_5316_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_Update/ca
      -- 
    ca_5953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2006_inst_ack_1, ack => convTransposeB_CP_5316_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	92 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109__exit__
      -- CP-element group 36: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/$exit
      -- CP-element group 36: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/$entry
      -- CP-element group 36: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2112/$entry
      -- CP-element group 36: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- 
    convTransposeB_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(33) & convTransposeB_CP_5316_elements(35);
      gj_convTransposeB_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	94 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_Sample/ra
      -- 
    ra_5965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2128_inst_ack_0, ack => convTransposeB_CP_5316_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	94 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_Sample/rr
      -- 
    ca_5970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2128_inst_ack_1, ack => convTransposeB_CP_5316_elements(38)); -- 
    rr_5978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(38), ack => type_cast_2158_inst_req_0); -- 
    rr_6088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(38), ack => type_cast_2189_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_Sample/ra
      -- 
    ra_5979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2158_inst_ack_0, ack => convTransposeB_CP_5316_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	94 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_Sample/req
      -- 
    ca_5984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2158_inst_ack_1, ack => convTransposeB_CP_5316_elements(40)); -- 
    req_6009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(40), ack => array_obj_ref_2164_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_Sample/ack
      -- 
    ack_6010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2164_index_offset_ack_0, ack => convTransposeB_CP_5316_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	94 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_request/req
      -- 
    ack_6015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2164_index_offset_ack_1, ack => convTransposeB_CP_5316_elements(42)); -- 
    req_6024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(42), ack => addr_of_2165_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_request/ack
      -- 
    ack_6025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2165_final_reg_ack_0, ack => convTransposeB_CP_5316_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	94 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Sample/word_access_start/word_0/rr
      -- 
    ack_6030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2165_final_reg_ack_1, ack => convTransposeB_CP_5316_elements(44)); -- 
    rr_6063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(44), ack => ptr_deref_2169_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Sample/word_access_start/word_0/ra
      -- 
    ra_6064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2169_load_0_ack_0, ack => convTransposeB_CP_5316_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	94 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/ptr_deref_2169_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/ptr_deref_2169_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/ptr_deref_2169_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/ptr_deref_2169_Merge/merge_ack
      -- 
    ca_6075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2169_load_0_ack_1, ack => convTransposeB_CP_5316_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_Sample/ra
      -- 
    ra_6089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_0, ack => convTransposeB_CP_5316_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	94 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_Sample/req
      -- 
    ca_6094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_1, ack => convTransposeB_CP_5316_elements(48)); -- 
    req_6119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(48), ack => array_obj_ref_2195_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_Sample/ack
      -- 
    ack_6120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2195_index_offset_ack_0, ack => convTransposeB_CP_5316_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	94 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_request/req
      -- 
    ack_6125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2195_index_offset_ack_1, ack => convTransposeB_CP_5316_elements(50)); -- 
    req_6134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(50), ack => addr_of_2196_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_request/ack
      -- 
    ack_6135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2196_final_reg_ack_0, ack => convTransposeB_CP_5316_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	94 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_word_addrgen/root_register_ack
      -- 
    ack_6140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2196_final_reg_ack_1, ack => convTransposeB_CP_5316_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/ptr_deref_2199_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/ptr_deref_2199_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/ptr_deref_2199_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/ptr_deref_2199_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/word_access_start/word_0/rr
      -- 
    rr_6178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(53), ack => ptr_deref_2199_store_0_req_0); -- 
    convTransposeB_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(46) & convTransposeB_CP_5316_elements(52);
      gj_convTransposeB_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Sample/word_access_start/word_0/ra
      -- 
    ra_6179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2199_store_0_ack_0, ack => convTransposeB_CP_5316_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	94 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Update/word_access_complete/word_0/ca
      -- 
    ca_6190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2199_store_0_ack_1, ack => convTransposeB_CP_5316_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	94 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_Sample/ra
      -- 
    ra_6199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2205_inst_ack_0, ack => convTransposeB_CP_5316_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	94 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_Update/ca
      -- 
    ca_6204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2205_inst_ack_1, ack => convTransposeB_CP_5316_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217__exit__
      -- CP-element group 58: 	 branch_block_stmt_1842/if_stmt_2218__entry__
      -- CP-element group 58: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/$exit
      -- CP-element group 58: 	 branch_block_stmt_1842/if_stmt_2218_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1842/if_stmt_2218_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_1842/if_stmt_2218_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_1842/if_stmt_2218_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_1842/R_cmp_2219_place
      -- CP-element group 58: 	 branch_block_stmt_1842/if_stmt_2218_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1842/if_stmt_2218_else_link/$entry
      -- 
    branch_req_6212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(58), ack => if_stmt_2218_branch_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(41) & convTransposeB_CP_5316_elements(49) & convTransposeB_CP_5316_elements(55) & convTransposeB_CP_5316_elements(57);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	89 
    -- CP-element group 59: 	90 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_1842/merge_stmt_2224_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_1842/merge_stmt_2224__exit__
      -- CP-element group 59: 	 branch_block_stmt_1842/assign_stmt_2230__entry__
      -- CP-element group 59: 	 branch_block_stmt_1842/assign_stmt_2230__exit__
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/merge_stmt_2224_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1842/merge_stmt_2224_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1842/merge_stmt_2224_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1842/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/if_stmt_2218_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1842/if_stmt_2218_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_1842/assign_stmt_2230/$entry
      -- CP-element group 59: 	 branch_block_stmt_1842/assign_stmt_2230/$exit
      -- 
    if_choice_transition_6217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2218_branch_ack_1, ack => convTransposeB_CP_5316_elements(59)); -- 
    cr_6445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(59), ack => type_cast_2115_inst_req_1); -- 
    rr_6440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(59), ack => type_cast_2115_inst_req_0); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (18) 
      -- CP-element group 60: 	 branch_block_stmt_1842/merge_stmt_2232_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_1842/merge_stmt_2232__exit__
      -- CP-element group 60: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248__entry__
      -- CP-element group 60: 	 branch_block_stmt_1842/merge_stmt_2232_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_1842/merge_stmt_2232_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_1842/merge_stmt_2232_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_1842/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1842/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_1842/if_stmt_2218_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_1842/if_stmt_2218_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_1842/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/$entry
      -- CP-element group 60: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_Update/cr
      -- 
    else_choice_transition_6221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2218_branch_ack_0, ack => convTransposeB_CP_5316_elements(60)); -- 
    rr_6237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(60), ack => type_cast_2242_inst_req_0); -- 
    cr_6242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(60), ack => type_cast_2242_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_Sample/ra
      -- 
    ra_6238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2242_inst_ack_0, ack => convTransposeB_CP_5316_elements(61)); -- 
    -- CP-element group 62:  branch  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248__exit__
      -- CP-element group 62: 	 branch_block_stmt_1842/if_stmt_2249__entry__
      -- CP-element group 62: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/$exit
      -- CP-element group 62: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1842/assign_stmt_2238_to_assign_stmt_2248/type_cast_2242_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1842/if_stmt_2249_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1842/if_stmt_2249_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_1842/if_stmt_2249_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_1842/if_stmt_2249_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_1842/R_cmp77_2250_place
      -- CP-element group 62: 	 branch_block_stmt_1842/if_stmt_2249_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1842/if_stmt_2249_else_link/$entry
      -- 
    ca_6243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2242_inst_ack_1, ack => convTransposeB_CP_5316_elements(62)); -- 
    branch_req_6251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(62), ack => if_stmt_2249_branch_req_0); -- 
    -- CP-element group 63:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (18) 
      -- CP-element group 63: 	 branch_block_stmt_1842/merge_stmt_2255_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_1842/merge_stmt_2255__exit__
      -- CP-element group 63: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271__entry__
      -- CP-element group 63: 	 branch_block_stmt_1842/merge_stmt_2255_PhiAck/dummy
      -- CP-element group 63: 	 branch_block_stmt_1842/merge_stmt_2255_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_1842/merge_stmt_2255_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_1842/ifx_xelse_ifx_xthen79_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1842/ifx_xelse_ifx_xthen79_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_1842/if_stmt_2249_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_1842/if_stmt_2249_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_1842/ifx_xelse_ifx_xthen79
      -- CP-element group 63: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/$entry
      -- CP-element group 63: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_Update/cr
      -- 
    if_choice_transition_6256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2249_branch_ack_1, ack => convTransposeB_CP_5316_elements(63)); -- 
    rr_6273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(63), ack => type_cast_2270_inst_req_0); -- 
    cr_6278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(63), ack => type_cast_2270_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	95 
    -- CP-element group 64: 	96 
    -- CP-element group 64: 	98 
    -- CP-element group 64: 	99 
    -- CP-element group 64:  members (20) 
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/$entry
      -- CP-element group 64: 	 branch_block_stmt_1842/if_stmt_2249_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1842/if_stmt_2249_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend
      -- 
    else_choice_transition_6260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2249_branch_ack_0, ack => convTransposeB_CP_5316_elements(64)); -- 
    rr_6514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(64), ack => type_cast_2279_inst_req_0); -- 
    cr_6519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(64), ack => type_cast_2279_inst_req_1); -- 
    cr_6542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(64), ack => type_cast_2285_inst_req_1); -- 
    rr_6537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(64), ack => type_cast_2285_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_Sample/ra
      -- 
    ra_6274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2270_inst_ack_0, ack => convTransposeB_CP_5316_elements(65)); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	103 
    -- CP-element group 66: 	105 
    -- CP-element group 66: 	106 
    -- CP-element group 66:  members (23) 
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271__exit__
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/$exit
      -- CP-element group 66: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1842/assign_stmt_2261_to_assign_stmt_2271/type_cast_2270_Update/ca
      -- 
    ca_6279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2270_inst_ack_1, ack => convTransposeB_CP_5316_elements(66)); -- 
    cr_6591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(66), ack => type_cast_2283_inst_req_1); -- 
    cr_6568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(66), ack => type_cast_2277_inst_req_1); -- 
    rr_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(66), ack => type_cast_2277_inst_req_0); -- 
    rr_6586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(66), ack => type_cast_2283_inst_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	112 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_Sample/ra
      -- 
    ra_6291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2290_inst_ack_0, ack => convTransposeB_CP_5316_elements(67)); -- 
    -- CP-element group 68:  branch  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	112 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (13) 
      -- CP-element group 68: 	 branch_block_stmt_1842/if_stmt_2297_else_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296__exit__
      -- CP-element group 68: 	 branch_block_stmt_1842/if_stmt_2297__entry__
      -- CP-element group 68: 	 branch_block_stmt_1842/if_stmt_2297_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1842/if_stmt_2297_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1842/if_stmt_2297_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1842/if_stmt_2297_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1842/R_cmp89_2298_place
      -- CP-element group 68: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/$exit
      -- CP-element group 68: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_1842/if_stmt_2297_dead_link/$entry
      -- 
    ca_6296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2290_inst_ack_1, ack => convTransposeB_CP_5316_elements(68)); -- 
    branch_req_6304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(68), ack => if_stmt_2297_branch_req_0); -- 
    -- CP-element group 69:  merge  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (15) 
      -- CP-element group 69: 	 branch_block_stmt_1842/if_stmt_2297_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1842/merge_stmt_2303_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1842/merge_stmt_2303__exit__
      -- CP-element group 69: 	 branch_block_stmt_1842/assign_stmt_2307__entry__
      -- CP-element group 69: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_Sample/req
      -- CP-element group 69: 	 branch_block_stmt_1842/if_stmt_2297_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1842/merge_stmt_2303_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1842/merge_stmt_2303_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1842/merge_stmt_2303_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1842/ifx_xend_whilex_xend
      -- CP-element group 69: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_1842/assign_stmt_2307/$entry
      -- CP-element group 69: 	 branch_block_stmt_1842/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1842/ifx_xend_whilex_xend_PhiReq/$entry
      -- 
    if_choice_transition_6309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2297_branch_ack_1, ack => convTransposeB_CP_5316_elements(69)); -- 
    req_6326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(69), ack => WPIPE_Block1_done_2305_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70: 	79 
    -- CP-element group 70: 	81 
    -- CP-element group 70: 	82 
    -- CP-element group 70:  members (20) 
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1842/if_stmt_2297_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1842/if_stmt_2297_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/$entry
      -- 
    else_choice_transition_6313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2297_branch_ack_0, ack => convTransposeB_CP_5316_elements(70)); -- 
    cr_6413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(70), ack => type_cast_1989_inst_req_1); -- 
    rr_6408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(70), ack => type_cast_1989_inst_req_0); -- 
    cr_6390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(70), ack => type_cast_1996_inst_req_1); -- 
    rr_6385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(70), ack => type_cast_1996_inst_req_0); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_Update/req
      -- CP-element group 71: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_sample_completed_
      -- 
    ack_6327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2305_inst_ack_0, ack => convTransposeB_CP_5316_elements(71)); -- 
    req_6331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(71), ack => WPIPE_Block1_done_2305_inst_req_1); -- 
    -- CP-element group 72:  transition  place  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (16) 
      -- CP-element group 72: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_Update/ack
      -- CP-element group 72: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1842/return___PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_1842/merge_stmt_2309_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1842/merge_stmt_2309_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_1842/merge_stmt_2309_PhiAck/$exit
      -- CP-element group 72: 	 $exit
      -- CP-element group 72: 	 branch_block_stmt_1842/$exit
      -- CP-element group 72: 	 branch_block_stmt_1842/branch_block_stmt_1842__exit__
      -- CP-element group 72: 	 branch_block_stmt_1842/merge_stmt_2309_PhiAck/dummy
      -- CP-element group 72: 	 branch_block_stmt_1842/assign_stmt_2307__exit__
      -- CP-element group 72: 	 branch_block_stmt_1842/return__
      -- CP-element group 72: 	 branch_block_stmt_1842/merge_stmt_2309__exit__
      -- CP-element group 72: 	 branch_block_stmt_1842/return___PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_1842/assign_stmt_2307/WPIPE_Block1_done_2305_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1842/assign_stmt_2307/$exit
      -- 
    ack_6332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2305_inst_ack_1, ack => convTransposeB_CP_5316_elements(72)); -- 
    -- CP-element group 73:  transition  output  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/$exit
      -- CP-element group 73: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_req
      -- CP-element group 73: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1994_konst_delay_trans
      -- CP-element group 73: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/$exit
      -- 
    phi_stmt_1990_req_6343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1990_req_6343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(73), ack => phi_stmt_1990_req_0); -- 
    -- Element group convTransposeB_CP_5316_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => convTransposeB_CP_5316_elements(31), ack => convTransposeB_CP_5316_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	31 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Sample/$exit
      -- 
    ra_6360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1987_inst_ack_0, ack => convTransposeB_CP_5316_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	31 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Update/ca
      -- 
    ca_6365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1987_inst_ack_1, ack => convTransposeB_CP_5316_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/$exit
      -- CP-element group 76: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_req
      -- CP-element group 76: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/$exit
      -- CP-element group 76: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/$exit
      -- 
    phi_stmt_1984_req_6366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1984_req_6366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(76), ack => phi_stmt_1984_req_0); -- 
    convTransposeB_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(74) & convTransposeB_CP_5316_elements(75);
      gj_convTransposeB_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	85 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1842/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(73) & convTransposeB_CP_5316_elements(76);
      gj_convTransposeB_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/Sample/$exit
      -- 
    ra_6386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1996_inst_ack_0, ack => convTransposeB_CP_5316_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	70 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/Update/ca
      -- CP-element group 79: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/Update/$exit
      -- 
    ca_6391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1996_inst_ack_1, ack => convTransposeB_CP_5316_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	84 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_req
      -- CP-element group 80: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/type_cast_1996/$exit
      -- CP-element group 80: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/phi_stmt_1990_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1990/$exit
      -- 
    phi_stmt_1990_req_6392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1990_req_6392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(80), ack => phi_stmt_1990_req_1); -- 
    convTransposeB_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(78) & convTransposeB_CP_5316_elements(79);
      gj_convTransposeB_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	70 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Sample/$exit
      -- 
    ra_6409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1989_inst_ack_0, ack => convTransposeB_CP_5316_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Update/ca
      -- 
    ca_6414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1989_inst_ack_1, ack => convTransposeB_CP_5316_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/$exit
      -- CP-element group 83: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/$exit
      -- CP-element group 83: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/$exit
      -- CP-element group 83: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1984/phi_stmt_1984_req
      -- 
    phi_stmt_1984_req_6415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1984_req_6415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(83), ack => phi_stmt_1984_req_1); -- 
    convTransposeB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(81) & convTransposeB_CP_5316_elements(82);
      gj_convTransposeB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1842/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(80) & convTransposeB_CP_5316_elements(83);
      gj_convTransposeB_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  merge  fork  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	77 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1842/merge_stmt_1983_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1842/merge_stmt_1983_PhiAck/$entry
      -- 
    convTransposeB_CP_5316_elements(85) <= OrReduce(convTransposeB_CP_5316_elements(77) & convTransposeB_CP_5316_elements(84));
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1842/merge_stmt_1983_PhiAck/phi_stmt_1984_ack
      -- 
    phi_stmt_1984_ack_6420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1984_ack_0, ack => convTransposeB_CP_5316_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1842/merge_stmt_1983_PhiAck/phi_stmt_1990_ack
      -- 
    phi_stmt_1990_ack_6421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1990_ack_0, ack => convTransposeB_CP_5316_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  place  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	32 
    -- CP-element group 88: 	33 
    -- CP-element group 88: 	34 
    -- CP-element group 88: 	35 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_1842/merge_stmt_1983__exit__
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109__entry__
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/$entry
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2001_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1842/assign_stmt_2002_to_assign_stmt_2109/type_cast_2006_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1842/merge_stmt_1983_PhiAck/$exit
      -- 
    rr_5933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(88), ack => type_cast_2001_inst_req_0); -- 
    cr_5938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(88), ack => type_cast_2001_inst_req_1); -- 
    rr_5947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(88), ack => type_cast_2006_inst_req_0); -- 
    cr_5952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(88), ack => type_cast_2006_inst_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(86) & convTransposeB_CP_5316_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	59 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/Sample/$exit
      -- 
    ra_6441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2115_inst_ack_0, ack => convTransposeB_CP_5316_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	59 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/Update/ca
      -- 
    ca_6446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2115_inst_ack_1, ack => convTransposeB_CP_5316_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2115/$exit
      -- CP-element group 91: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/$exit
      -- CP-element group 91: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 91: 	 branch_block_stmt_1842/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_req
      -- 
    phi_stmt_2112_req_6447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2112_req_6447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(91), ack => phi_stmt_2112_req_0); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(89) & convTransposeB_CP_5316_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  output  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	36 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_req
      -- CP-element group 92: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/type_cast_2118_konst_delay_trans
      -- CP-element group 92: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2112/phi_stmt_2112_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2112/$exit
      -- CP-element group 92: 	 branch_block_stmt_1842/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_2112_req_6458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2112_req_6458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(92), ack => phi_stmt_2112_req_1); -- 
    -- Element group convTransposeB_CP_5316_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => convTransposeB_CP_5316_elements(36), ack => convTransposeB_CP_5316_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  merge  transition  place  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1842/merge_stmt_2111_PhiReqMerge
      -- CP-element group 93: 	 branch_block_stmt_1842/merge_stmt_2111_PhiAck/$entry
      -- 
    convTransposeB_CP_5316_elements(93) <= OrReduce(convTransposeB_CP_5316_elements(91) & convTransposeB_CP_5316_elements(92));
    -- CP-element group 94:  fork  transition  place  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	40 
    -- CP-element group 94: 	46 
    -- CP-element group 94: 	42 
    -- CP-element group 94: 	48 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	38 
    -- CP-element group 94: 	44 
    -- CP-element group 94: 	50 
    -- CP-element group 94: 	52 
    -- CP-element group 94: 	55 
    -- CP-element group 94: 	56 
    -- CP-element group 94: 	57 
    -- CP-element group 94:  members (45) 
      -- CP-element group 94: 	 branch_block_stmt_1842/merge_stmt_2111__exit__
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217__entry__
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2128_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2158_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2164_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2165_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2169_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2189_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/array_obj_ref_2195_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1842/merge_stmt_2111_PhiAck/phi_stmt_2112_ack
      -- CP-element group 94: 	 branch_block_stmt_1842/merge_stmt_2111_PhiAck/$exit
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/addr_of_2196_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/ptr_deref_2199_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1842/assign_stmt_2125_to_assign_stmt_2217/type_cast_2205_Update/cr
      -- 
    phi_stmt_2112_ack_6463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2112_ack_0, ack => convTransposeB_CP_5316_elements(94)); -- 
    rr_5964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => type_cast_2128_inst_req_0); -- 
    cr_5969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => type_cast_2128_inst_req_1); -- 
    cr_5983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => type_cast_2158_inst_req_1); -- 
    req_6014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => array_obj_ref_2164_index_offset_req_1); -- 
    req_6029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => addr_of_2165_final_reg_req_1); -- 
    cr_6074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => ptr_deref_2169_load_0_req_1); -- 
    cr_6093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => type_cast_2189_inst_req_1); -- 
    req_6124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => array_obj_ref_2195_index_offset_req_1); -- 
    req_6139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => addr_of_2196_final_reg_req_1); -- 
    cr_6189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => ptr_deref_2199_store_0_req_1); -- 
    rr_6198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => type_cast_2205_inst_req_0); -- 
    cr_6203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(94), ack => type_cast_2205_inst_req_1); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	64 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/Sample/ra
      -- 
    ra_6515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2279_inst_ack_0, ack => convTransposeB_CP_5316_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	64 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/Update/ca
      -- 
    ca_6520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2279_inst_ack_1, ack => convTransposeB_CP_5316_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/$exit
      -- CP-element group 97: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/$exit
      -- CP-element group 97: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2279/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_req
      -- 
    phi_stmt_2274_req_6521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2274_req_6521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(97), ack => phi_stmt_2274_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(95) & convTransposeB_CP_5316_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	64 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/Sample/$exit
      -- 
    ra_6538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2285_inst_ack_0, ack => convTransposeB_CP_5316_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	64 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/Update/ca
      -- CP-element group 99: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/Update/$exit
      -- 
    ca_6543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2285_inst_ack_1, ack => convTransposeB_CP_5316_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/$exit
      -- CP-element group 100: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_req
      -- CP-element group 100: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2285/$exit
      -- CP-element group 100: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/$exit
      -- 
    phi_stmt_2280_req_6544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2280_req_6544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(100), ack => phi_stmt_2280_req_1); -- 
    convTransposeB_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(98) & convTransposeB_CP_5316_elements(99);
      gj_convTransposeB_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	109 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1842/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(97) & convTransposeB_CP_5316_elements(100);
      gj_convTransposeB_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/Sample/$exit
      -- 
    ra_6564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2277_inst_ack_0, ack => convTransposeB_CP_5316_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/Update/ca
      -- CP-element group 103: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/Update/$exit
      -- 
    ca_6569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2277_inst_ack_1, ack => convTransposeB_CP_5316_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_req
      -- CP-element group 104: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/type_cast_2277/$exit
      -- CP-element group 104: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/phi_stmt_2274_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2274/$exit
      -- 
    phi_stmt_2274_req_6570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2274_req_6570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(104), ack => phi_stmt_2274_req_0); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(102) & convTransposeB_CP_5316_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	66 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/Sample/ra
      -- 
    ra_6587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2283_inst_ack_0, ack => convTransposeB_CP_5316_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	66 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/Update/$exit
      -- 
    ca_6592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2283_inst_ack_1, ack => convTransposeB_CP_5316_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/$exit
      -- CP-element group 107: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_req
      -- CP-element group 107: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/type_cast_2283/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/phi_stmt_2280_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2280/$exit
      -- 
    phi_stmt_2280_req_6593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2280_req_6593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(107), ack => phi_stmt_2280_req_0); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(105) & convTransposeB_CP_5316_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1842/ifx_xthen79_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(104) & convTransposeB_CP_5316_elements(107);
      gj_convTransposeB_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	101 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1842/merge_stmt_2273_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_1842/merge_stmt_2273_PhiAck/$entry
      -- 
    convTransposeB_CP_5316_elements(109) <= OrReduce(convTransposeB_CP_5316_elements(101) & convTransposeB_CP_5316_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1842/merge_stmt_2273_PhiAck/phi_stmt_2274_ack
      -- 
    phi_stmt_2274_ack_6598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2274_ack_0, ack => convTransposeB_CP_5316_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1842/merge_stmt_2273_PhiAck/phi_stmt_2280_ack
      -- 
    phi_stmt_2280_ack_6599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2280_ack_0, ack => convTransposeB_CP_5316_elements(111)); -- 
    -- CP-element group 112:  join  fork  transition  place  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: 	68 
    -- CP-element group 112:  members (10) 
      -- CP-element group 112: 	 branch_block_stmt_1842/merge_stmt_2273_PhiAck/$exit
      -- CP-element group 112: 	 branch_block_stmt_1842/merge_stmt_2273__exit__
      -- CP-element group 112: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296__entry__
      -- CP-element group 112: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/$entry
      -- CP-element group 112: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1842/assign_stmt_2291_to_assign_stmt_2296/type_cast_2290_Update/cr
      -- 
    rr_6290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(112), ack => type_cast_2290_inst_req_0); -- 
    cr_6295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5316_elements(112), ack => type_cast_2290_inst_req_1); -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5316_elements(110) & convTransposeB_CP_5316_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5316_elements(112), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2071_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2092_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2152_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2183_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1908_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1908_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom61_2194_resized : std_logic_vector(13 downto 0);
    signal R_idxprom61_2194_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2163_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2163_scaled : std_logic_vector(13 downto 0);
    signal add17_2134 : std_logic_vector(31 downto 0);
    signal add25_2032 : std_logic_vector(31 downto 0);
    signal add36_2047 : std_logic_vector(31 downto 0);
    signal add51_2104 : std_logic_vector(31 downto 0);
    signal add53_2139 : std_logic_vector(31 downto 0);
    signal add66_2212 : std_logic_vector(31 downto 0);
    signal add_2017 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2164_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2164_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2164_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2164_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2164_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2164_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2195_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2195_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2195_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2195_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2195_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2195_root_address : std_logic_vector(13 downto 0);
    signal arrayidx62_2197 : std_logic_vector(31 downto 0);
    signal arrayidx_2166 : std_logic_vector(31 downto 0);
    signal call_1845 : std_logic_vector(15 downto 0);
    signal cmp77_2248 : std_logic_vector(0 downto 0);
    signal cmp89_2296 : std_logic_vector(0 downto 0);
    signal cmp_2217 : std_logic_vector(0 downto 0);
    signal conv12_2002 : std_logic_vector(31 downto 0);
    signal conv15_2007 : std_logic_vector(31 downto 0);
    signal conv22_1894 : std_logic_vector(31 downto 0);
    signal conv27_1913 : std_logic_vector(31 downto 0);
    signal conv33_1927 : std_logic_vector(31 downto 0);
    signal conv46_2073 : std_logic_vector(31 downto 0);
    signal conv49_2094 : std_logic_vector(31 downto 0);
    signal conv65_2206 : std_logic_vector(31 downto 0);
    signal conv75_2243 : std_logic_vector(31 downto 0);
    signal conv84_2271 : std_logic_vector(15 downto 0);
    signal conv86_2291 : std_logic_vector(31 downto 0);
    signal conv9102_2129 : std_logic_vector(31 downto 0);
    signal conv_1868 : std_logic_vector(15 downto 0);
    signal div83_2267 : std_logic_vector(31 downto 0);
    signal div88_1981 : std_logic_vector(31 downto 0);
    signal div_1864 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1971 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1854 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1876 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1886 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1902 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1919 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1935 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1947 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1959 : std_logic_vector(31 downto 0);
    signal idxprom61_2190 : std_logic_vector(63 downto 0);
    signal idxprom_2159 : std_logic_vector(63 downto 0);
    signal inc81_2261 : std_logic_vector(15 downto 0);
    signal inc_2238 : std_logic_vector(15 downto 0);
    signal indvar_2112 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2230 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2280 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1990 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1984 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2274 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2125 : std_logic_vector(15 downto 0);
    signal mul16_2022 : std_logic_vector(31 downto 0);
    signal mul23_2027 : std_logic_vector(31 downto 0);
    signal mul34_2042 : std_logic_vector(31 downto 0);
    signal mul50_2099 : std_logic_vector(31 downto 0);
    signal mul52_2109 : std_logic_vector(31 downto 0);
    signal mul_2012 : std_logic_vector(31 downto 0);
    signal ptr_deref_1857_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1857_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1857_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1857_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1857_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1879_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1879_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1879_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1879_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1879_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1889_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1889_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1889_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1889_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1889_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1905_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1905_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1905_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1905_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1905_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1922_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1922_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1922_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1922_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1922_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1938_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1938_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1938_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1938_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1938_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1950_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1950_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1950_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1950_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1950_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1962_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1962_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1962_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1962_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1962_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1974_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1974_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1974_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1974_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1974_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2169_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2169_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2199_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2199_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2199_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2199_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2199_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2199_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext103_2085 : std_logic_vector(31 downto 0);
    signal sext105_2145 : std_logic_vector(31 downto 0);
    signal sext106_2176 : std_logic_vector(31 downto 0);
    signal sext_2064 : std_logic_vector(31 downto 0);
    signal shr60_2185 : std_logic_vector(31 downto 0);
    signal shr_2154 : std_logic_vector(31 downto 0);
    signal sub28_2079 : std_logic_vector(31 downto 0);
    signal sub39_2052 : std_logic_vector(31 downto 0);
    signal sub40_2058 : std_logic_vector(31 downto 0);
    signal sub_2037 : std_logic_vector(31 downto 0);
    signal tmp10_1880 : std_logic_vector(31 downto 0);
    signal tmp21_1890 : std_logic_vector(15 downto 0);
    signal tmp24_1906 : std_logic_vector(31 downto 0);
    signal tmp26_1909 : std_logic_vector(15 downto 0);
    signal tmp32_1923 : std_logic_vector(15 downto 0);
    signal tmp35_1939 : std_logic_vector(31 downto 0);
    signal tmp44_1951 : std_logic_vector(31 downto 0);
    signal tmp47_1963 : std_logic_vector(31 downto 0);
    signal tmp57_2170 : std_logic_vector(63 downto 0);
    signal tmp87_1975 : std_logic_vector(31 downto 0);
    signal tmp_1858 : std_logic_vector(31 downto 0);
    signal type_cast_1862_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1979_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1987_wire : std_logic_vector(15 downto 0);
    signal type_cast_1989_wire : std_logic_vector(15 downto 0);
    signal type_cast_1994_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1996_wire : std_logic_vector(15 downto 0);
    signal type_cast_2000_wire : std_logic_vector(31 downto 0);
    signal type_cast_2005_wire : std_logic_vector(31 downto 0);
    signal type_cast_2056_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2062_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2067_wire : std_logic_vector(31 downto 0);
    signal type_cast_2070_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2077_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2083_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2088_wire : std_logic_vector(31 downto 0);
    signal type_cast_2091_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2115_wire : std_logic_vector(15 downto 0);
    signal type_cast_2118_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2123_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2143_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2148_wire : std_logic_vector(31 downto 0);
    signal type_cast_2151_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2157_wire : std_logic_vector(63 downto 0);
    signal type_cast_2174_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2179_wire : std_logic_vector(31 downto 0);
    signal type_cast_2182_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2188_wire : std_logic_vector(63 downto 0);
    signal type_cast_2204_wire : std_logic_vector(31 downto 0);
    signal type_cast_2210_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2228_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2236_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2241_wire : std_logic_vector(31 downto 0);
    signal type_cast_2259_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2265_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2277_wire : std_logic_vector(15 downto 0);
    signal type_cast_2279_wire : std_logic_vector(15 downto 0);
    signal type_cast_2283_wire : std_logic_vector(15 downto 0);
    signal type_cast_2285_wire : std_logic_vector(15 downto 0);
    signal type_cast_2289_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1908_word_address_0 <= "0";
    array_obj_ref_2164_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2164_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2164_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2164_resized_base_address <= "00000000000000";
    array_obj_ref_2195_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2195_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2195_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2195_resized_base_address <= "00000000000000";
    iNsTr_10_1971 <= "00000000000000000000000000000010";
    iNsTr_2_1854 <= "00000000000000000000000000000011";
    iNsTr_3_1876 <= "00000000000000000000000000000100";
    iNsTr_4_1886 <= "00000000000000000000000000000000";
    iNsTr_5_1902 <= "00000000000000000000000000000011";
    iNsTr_6_1919 <= "00000000000000000000000000000001";
    iNsTr_7_1935 <= "00000000000000000000000000000100";
    iNsTr_8_1947 <= "00000000000000000000000000000100";
    iNsTr_9_1959 <= "00000000000000000000000000000011";
    ptr_deref_1857_word_offset_0 <= "0000000";
    ptr_deref_1879_word_offset_0 <= "0000000";
    ptr_deref_1889_word_offset_0 <= "0";
    ptr_deref_1905_word_offset_0 <= "0000000";
    ptr_deref_1922_word_offset_0 <= "0";
    ptr_deref_1938_word_offset_0 <= "0000000";
    ptr_deref_1950_word_offset_0 <= "0000000";
    ptr_deref_1962_word_offset_0 <= "0000000";
    ptr_deref_1974_word_offset_0 <= "0000000";
    ptr_deref_2169_word_offset_0 <= "00000000000000";
    ptr_deref_2199_word_offset_0 <= "00000000000000";
    type_cast_1862_wire_constant <= "00000000000000000000000000000001";
    type_cast_1979_wire_constant <= "00000000000000000000000000000001";
    type_cast_1994_wire_constant <= "0000000000000000";
    type_cast_2056_wire_constant <= "00000000000000000000000000010000";
    type_cast_2062_wire_constant <= "11111111111111110000000000000000";
    type_cast_2070_wire_constant <= "00000000000000000000000000010000";
    type_cast_2077_wire_constant <= "00000000000000000000000000010000";
    type_cast_2083_wire_constant <= "11111111111111110000000000000000";
    type_cast_2091_wire_constant <= "00000000000000000000000000010000";
    type_cast_2118_wire_constant <= "0000000000000000";
    type_cast_2123_wire_constant <= "0000000000000100";
    type_cast_2143_wire_constant <= "00000000000000000000000000010000";
    type_cast_2151_wire_constant <= "00000000000000000000000000010010";
    type_cast_2174_wire_constant <= "00000000000000000000000000010000";
    type_cast_2182_wire_constant <= "00000000000000000000000000010010";
    type_cast_2210_wire_constant <= "00000000000000000000000000000100";
    type_cast_2228_wire_constant <= "0000000000000001";
    type_cast_2236_wire_constant <= "0000000000000001";
    type_cast_2259_wire_constant <= "0000000000000001";
    type_cast_2265_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1984: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1987_wire & type_cast_1989_wire;
      req <= phi_stmt_1984_req_0 & phi_stmt_1984_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1984",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1984_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1984,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1984
    phi_stmt_1990: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1994_wire_constant & type_cast_1996_wire;
      req <= phi_stmt_1990_req_0 & phi_stmt_1990_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1990",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1990_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1990,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1990
    phi_stmt_2112: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2115_wire & type_cast_2118_wire_constant;
      req <= phi_stmt_2112_req_0 & phi_stmt_2112_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2112",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2112_ack_0,
          idata => idata,
          odata => indvar_2112,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2112
    phi_stmt_2274: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2277_wire & type_cast_2279_wire;
      req <= phi_stmt_2274_req_0 & phi_stmt_2274_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2274",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2274_ack_0,
          idata => idata,
          odata => input_dim1x_x2_2274,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2274
    phi_stmt_2280: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2283_wire & type_cast_2285_wire;
      req <= phi_stmt_2280_req_0 & phi_stmt_2280_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2280",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2280_ack_0,
          idata => idata,
          odata => input_dim0x_x0_2280,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2280
    addr_of_2165_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2165_final_reg_req_0;
      addr_of_2165_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2165_final_reg_req_1;
      addr_of_2165_final_reg_ack_1<= rack(0);
      addr_of_2165_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2165_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2164_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2166,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2196_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2196_final_reg_req_0;
      addr_of_2196_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2196_final_reg_req_1;
      addr_of_2196_final_reg_ack_1<= rack(0);
      addr_of_2196_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2196_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2195_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx62_2197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1867_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1867_inst_req_0;
      type_cast_1867_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1867_inst_req_1;
      type_cast_1867_inst_ack_1<= rack(0);
      type_cast_1867_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1867_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1864,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1868,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1893_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1893_inst_req_0;
      type_cast_1893_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1893_inst_req_1;
      type_cast_1893_inst_ack_1<= rack(0);
      type_cast_1893_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1893_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp21_1890,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1894,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1912_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1912_inst_req_0;
      type_cast_1912_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1912_inst_req_1;
      type_cast_1912_inst_ack_1<= rack(0);
      type_cast_1912_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1912_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26_1909,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_1913,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1926_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1926_inst_req_0;
      type_cast_1926_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1926_inst_req_1;
      type_cast_1926_inst_ack_1<= rack(0);
      type_cast_1926_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1926_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp32_1923,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1927,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1987_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1987_inst_req_0;
      type_cast_1987_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1987_inst_req_1;
      type_cast_1987_inst_ack_1<= rack(0);
      type_cast_1987_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1987_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_1868,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1987_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1989_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1989_inst_req_0;
      type_cast_1989_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1989_inst_req_1;
      type_cast_1989_inst_ack_1<= rack(0);
      type_cast_1989_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1989_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2274,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1989_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1996_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1996_inst_req_0;
      type_cast_1996_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1996_inst_req_1;
      type_cast_1996_inst_ack_1<= rack(0);
      type_cast_1996_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1996_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1996_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2001_inst_req_0;
      type_cast_2001_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2001_inst_req_1;
      type_cast_2001_inst_ack_1<= rack(0);
      type_cast_2001_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2000_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_2002,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2006_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2006_inst_req_0;
      type_cast_2006_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2006_inst_req_1;
      type_cast_2006_inst_ack_1<= rack(0);
      type_cast_2006_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2006_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2005_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_2007,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2067_inst
    process(sext_2064) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2064(31 downto 0);
      type_cast_2067_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2072_inst
    process(ASHR_i32_i32_2071_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2071_wire(31 downto 0);
      conv46_2073 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2088_inst
    process(sext103_2085) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2085(31 downto 0);
      type_cast_2088_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2093_inst
    process(ASHR_i32_i32_2092_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2092_wire(31 downto 0);
      conv49_2094 <= tmp_var; -- 
    end process;
    type_cast_2115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2115_inst_req_0;
      type_cast_2115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2115_inst_req_1;
      type_cast_2115_inst_ack_1<= rack(0);
      type_cast_2115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2115_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2128_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2128_inst_req_0;
      type_cast_2128_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2128_inst_req_1;
      type_cast_2128_inst_ack_1<= rack(0);
      type_cast_2128_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2128_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9102_2129,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2148_inst
    process(sext105_2145) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext105_2145(31 downto 0);
      type_cast_2148_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2153_inst
    process(ASHR_i32_i32_2152_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2152_wire(31 downto 0);
      shr_2154 <= tmp_var; -- 
    end process;
    type_cast_2158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2158_inst_req_0;
      type_cast_2158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2158_inst_req_1;
      type_cast_2158_inst_ack_1<= rack(0);
      type_cast_2158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2157_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2179_inst
    process(sext106_2176) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2176(31 downto 0);
      type_cast_2179_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2184_inst
    process(ASHR_i32_i32_2183_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2183_wire(31 downto 0);
      shr60_2185 <= tmp_var; -- 
    end process;
    type_cast_2189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2189_inst_req_0;
      type_cast_2189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2189_inst_req_1;
      type_cast_2189_inst_ack_1<= rack(0);
      type_cast_2189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2188_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom61_2190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2205_inst_req_0;
      type_cast_2205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2205_inst_req_1;
      type_cast_2205_inst_ack_1<= rack(0);
      type_cast_2205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2204_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2242_inst_req_0;
      type_cast_2242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2242_inst_req_1;
      type_cast_2242_inst_ack_1<= rack(0);
      type_cast_2242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2242_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2241_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2270_inst_req_0;
      type_cast_2270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2270_inst_req_1;
      type_cast_2270_inst_ack_1<= rack(0);
      type_cast_2270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div83_2267,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2277_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2277_inst_req_0;
      type_cast_2277_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2277_inst_req_1;
      type_cast_2277_inst_ack_1<= rack(0);
      type_cast_2277_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2277_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv84_2271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2277_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2279_inst_req_0;
      type_cast_2279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2279_inst_req_1;
      type_cast_2279_inst_ack_1<= rack(0);
      type_cast_2279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2279_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2283_inst_req_0;
      type_cast_2283_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2283_inst_req_1;
      type_cast_2283_inst_ack_1<= rack(0);
      type_cast_2283_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2283_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc81_2261,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2283_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2285_inst_req_0;
      type_cast_2285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2285_inst_req_1;
      type_cast_2285_inst_ack_1<= rack(0);
      type_cast_2285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_1990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2285_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2290_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2290_inst_req_0;
      type_cast_2290_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2290_inst_req_1;
      type_cast_2290_inst_ack_1<= rack(0);
      type_cast_2290_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2290_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2289_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2291,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1908_gather_scatter
    process(LOAD_padding_1908_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1908_data_0;
      ov(15 downto 0) := iv;
      tmp26_1909 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2164_index_1_rename
    process(R_idxprom_2163_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2163_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2163_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2164_index_1_resize
    process(idxprom_2159) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2159;
      ov := iv(13 downto 0);
      R_idxprom_2163_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2164_root_address_inst
    process(array_obj_ref_2164_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2164_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2164_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2195_index_1_rename
    process(R_idxprom61_2194_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom61_2194_resized;
      ov(13 downto 0) := iv;
      R_idxprom61_2194_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2195_index_1_resize
    process(idxprom61_2190) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom61_2190;
      ov := iv(13 downto 0);
      R_idxprom61_2194_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2195_root_address_inst
    process(array_obj_ref_2195_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2195_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2195_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1857_addr_0
    process(ptr_deref_1857_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1857_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1857_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1857_base_resize
    process(iNsTr_2_1854) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1854;
      ov := iv(6 downto 0);
      ptr_deref_1857_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1857_gather_scatter
    process(ptr_deref_1857_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1857_data_0;
      ov(31 downto 0) := iv;
      tmp_1858 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1857_root_address_inst
    process(ptr_deref_1857_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1857_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1857_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1879_addr_0
    process(ptr_deref_1879_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1879_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1879_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1879_base_resize
    process(iNsTr_3_1876) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1876;
      ov := iv(6 downto 0);
      ptr_deref_1879_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1879_gather_scatter
    process(ptr_deref_1879_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1879_data_0;
      ov(31 downto 0) := iv;
      tmp10_1880 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1879_root_address_inst
    process(ptr_deref_1879_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1879_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1879_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1889_addr_0
    process(ptr_deref_1889_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1889_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1889_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1889_base_resize
    process(iNsTr_4_1886) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1886;
      ov := iv(0 downto 0);
      ptr_deref_1889_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1889_gather_scatter
    process(ptr_deref_1889_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1889_data_0;
      ov(15 downto 0) := iv;
      tmp21_1890 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1889_root_address_inst
    process(ptr_deref_1889_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1889_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1889_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_addr_0
    process(ptr_deref_1905_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1905_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_base_resize
    process(iNsTr_5_1902) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1902;
      ov := iv(6 downto 0);
      ptr_deref_1905_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_gather_scatter
    process(ptr_deref_1905_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_data_0;
      ov(31 downto 0) := iv;
      tmp24_1906 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_root_address_inst
    process(ptr_deref_1905_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1905_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1922_addr_0
    process(ptr_deref_1922_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1922_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1922_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1922_base_resize
    process(iNsTr_6_1919) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1919;
      ov := iv(0 downto 0);
      ptr_deref_1922_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1922_gather_scatter
    process(ptr_deref_1922_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1922_data_0;
      ov(15 downto 0) := iv;
      tmp32_1923 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1922_root_address_inst
    process(ptr_deref_1922_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1922_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1922_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1938_addr_0
    process(ptr_deref_1938_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1938_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1938_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1938_base_resize
    process(iNsTr_7_1935) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1935;
      ov := iv(6 downto 0);
      ptr_deref_1938_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1938_gather_scatter
    process(ptr_deref_1938_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1938_data_0;
      ov(31 downto 0) := iv;
      tmp35_1939 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1938_root_address_inst
    process(ptr_deref_1938_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1938_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1938_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1950_addr_0
    process(ptr_deref_1950_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1950_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1950_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1950_base_resize
    process(iNsTr_8_1947) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1947;
      ov := iv(6 downto 0);
      ptr_deref_1950_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1950_gather_scatter
    process(ptr_deref_1950_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1950_data_0;
      ov(31 downto 0) := iv;
      tmp44_1951 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1950_root_address_inst
    process(ptr_deref_1950_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1950_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1950_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1962_addr_0
    process(ptr_deref_1962_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1962_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1962_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1962_base_resize
    process(iNsTr_9_1959) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1959;
      ov := iv(6 downto 0);
      ptr_deref_1962_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1962_gather_scatter
    process(ptr_deref_1962_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1962_data_0;
      ov(31 downto 0) := iv;
      tmp47_1963 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1962_root_address_inst
    process(ptr_deref_1962_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1962_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1962_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1974_addr_0
    process(ptr_deref_1974_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1974_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1974_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1974_base_resize
    process(iNsTr_10_1971) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1971;
      ov := iv(6 downto 0);
      ptr_deref_1974_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1974_gather_scatter
    process(ptr_deref_1974_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1974_data_0;
      ov(31 downto 0) := iv;
      tmp87_1975 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1974_root_address_inst
    process(ptr_deref_1974_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1974_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1974_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_addr_0
    process(ptr_deref_2169_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2169_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2169_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_base_resize
    process(arrayidx_2166) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2166;
      ov := iv(13 downto 0);
      ptr_deref_2169_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_gather_scatter
    process(ptr_deref_2169_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2169_data_0;
      ov(63 downto 0) := iv;
      tmp57_2170 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_root_address_inst
    process(ptr_deref_2169_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2169_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2169_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2199_addr_0
    process(ptr_deref_2199_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2199_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2199_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2199_base_resize
    process(arrayidx62_2197) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx62_2197;
      ov := iv(13 downto 0);
      ptr_deref_2199_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2199_gather_scatter
    process(tmp57_2170) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp57_2170;
      ov(63 downto 0) := iv;
      ptr_deref_2199_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2199_root_address_inst
    process(ptr_deref_2199_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2199_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2199_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2218_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2217;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2218_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2218_branch_req_0,
          ack0 => if_stmt_2218_branch_ack_0,
          ack1 => if_stmt_2218_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2249_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_2248;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2249_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2249_branch_req_0,
          ack0 => if_stmt_2249_branch_ack_0,
          ack1 => if_stmt_2249_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2297_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp89_2296;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2297_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2297_branch_req_0,
          ack0 => if_stmt_2297_branch_ack_0,
          ack1 => if_stmt_2297_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2229_inst
    process(indvar_2112) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2112, type_cast_2228_wire_constant, tmp_var);
      indvarx_xnext_2230 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2237_inst
    process(input_dim1x_x1x_xph_1984) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1984, type_cast_2236_wire_constant, tmp_var);
      inc_2238 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2260_inst
    process(input_dim0x_x2x_xph_1990) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_1990, type_cast_2259_wire_constant, tmp_var);
      inc81_2261 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2016_inst
    process(mul_2012, conv12_2002) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2012, conv12_2002, tmp_var);
      add_2017 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2031_inst
    process(mul23_2027, tmp24_1906) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul23_2027, tmp24_1906, tmp_var);
      add25_2032 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2046_inst
    process(mul34_2042, tmp35_1939) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul34_2042, tmp35_1939, tmp_var);
      add36_2047 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2063_inst
    process(sub40_2058) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub40_2058, type_cast_2062_wire_constant, tmp_var);
      sext_2064 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2084_inst
    process(sub28_2079) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub28_2079, type_cast_2083_wire_constant, tmp_var);
      sext103_2085 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2103_inst
    process(conv46_2073, mul50_2099) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv46_2073, mul50_2099, tmp_var);
      add51_2104 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2133_inst
    process(mul16_2022, conv9102_2129) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul16_2022, conv9102_2129, tmp_var);
      add17_2134 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2138_inst
    process(mul52_2109, conv9102_2129) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul52_2109, conv9102_2129, tmp_var);
      add53_2139 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2211_inst
    process(conv65_2206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv65_2206, type_cast_2210_wire_constant, tmp_var);
      add66_2212 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2071_inst
    process(type_cast_2067_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2067_wire, type_cast_2070_wire_constant, tmp_var);
      ASHR_i32_i32_2071_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2092_inst
    process(type_cast_2088_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2088_wire, type_cast_2091_wire_constant, tmp_var);
      ASHR_i32_i32_2092_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2152_inst
    process(type_cast_2148_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2148_wire, type_cast_2151_wire_constant, tmp_var);
      ASHR_i32_i32_2152_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2183_inst
    process(type_cast_2179_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2179_wire, type_cast_2182_wire_constant, tmp_var);
      ASHR_i32_i32_2183_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2247_inst
    process(conv75_2243, tmp_1858) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv75_2243, tmp_1858, tmp_var);
      cmp77_2248 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2295_inst
    process(conv86_2291, div88_1981) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv86_2291, div88_1981, tmp_var);
      cmp89_2296 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1863_inst
    process(tmp_1858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1858, type_cast_1862_wire_constant, tmp_var);
      div_1864 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1980_inst
    process(tmp87_1975) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp87_1975, type_cast_1979_wire_constant, tmp_var);
      div88_1981 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2266_inst
    process(tmp_1858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1858, type_cast_2265_wire_constant, tmp_var);
      div83_2267 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2124_inst
    process(indvar_2112) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2112, type_cast_2123_wire_constant, tmp_var);
      input_dim2x_x1_2125 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2011_inst
    process(tmp_1858, conv15_2007) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1858, conv15_2007, tmp_var);
      mul_2012 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2021_inst
    process(add_2017, tmp10_1880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2017, tmp10_1880, tmp_var);
      mul16_2022 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2026_inst
    process(conv22_1894, conv15_2007) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv22_1894, conv15_2007, tmp_var);
      mul23_2027 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2041_inst
    process(conv33_1927, conv12_2002) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_1927, conv12_2002, tmp_var);
      mul34_2042 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2098_inst
    process(tmp47_1963, conv49_2094) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp47_1963, conv49_2094, tmp_var);
      mul50_2099 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2108_inst
    process(add51_2104, tmp44_1951) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add51_2104, tmp44_1951, tmp_var);
      mul52_2109 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2057_inst
    process(sub39_2052) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub39_2052, type_cast_2056_wire_constant, tmp_var);
      sub40_2058 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2078_inst
    process(sub_2037) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2037, type_cast_2077_wire_constant, tmp_var);
      sub28_2079 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2144_inst
    process(add17_2134) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add17_2134, type_cast_2143_wire_constant, tmp_var);
      sext105_2145 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2175_inst
    process(add53_2139) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add53_2139, type_cast_2174_wire_constant, tmp_var);
      sext106_2176 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2036_inst
    process(add25_2032, conv27_1913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add25_2032, conv27_1913, tmp_var);
      sub_2037 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2051_inst
    process(add36_2047, conv27_1913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add36_2047, conv27_1913, tmp_var);
      sub39_2052 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2216_inst
    process(add66_2212, tmp10_1880) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add66_2212, tmp10_1880, tmp_var);
      cmp_2217 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_2164_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2163_scaled;
      array_obj_ref_2164_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2164_index_offset_req_0;
      array_obj_ref_2164_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2164_index_offset_req_1;
      array_obj_ref_2164_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_2195_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom61_2194_scaled;
      array_obj_ref_2195_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2195_index_offset_req_0;
      array_obj_ref_2195_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2195_index_offset_req_1;
      array_obj_ref_2195_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_2000_inst
    process(input_dim1x_x1x_xph_1984) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1984, tmp_var);
      type_cast_2000_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2005_inst
    process(input_dim0x_x2x_xph_1990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1990, tmp_var);
      type_cast_2005_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2157_inst
    process(shr_2154) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2154, tmp_var);
      type_cast_2157_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2188_inst
    process(shr60_2185) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr60_2185, tmp_var);
      type_cast_2188_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2204_inst
    process(input_dim2x_x1_2125) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2125, tmp_var);
      type_cast_2204_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2241_inst
    process(inc_2238) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2238, tmp_var);
      type_cast_2241_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2289_inst
    process(input_dim0x_x0_2280) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2280, tmp_var);
      type_cast_2289_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1908_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1908_load_0_req_0;
      LOAD_padding_1908_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1908_load_0_req_1;
      LOAD_padding_1908_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1908_word_address_0;
      LOAD_padding_1908_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1857_load_0 ptr_deref_1879_load_0 ptr_deref_1974_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1857_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1879_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1974_load_0_req_0;
      ptr_deref_1857_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1879_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1974_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1857_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1879_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1974_load_0_req_1;
      ptr_deref_1857_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1879_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1974_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1857_word_address_0 & ptr_deref_1879_word_address_0 & ptr_deref_1974_word_address_0;
      ptr_deref_1857_data_0 <= data_out(95 downto 64);
      ptr_deref_1879_data_0 <= data_out(63 downto 32);
      ptr_deref_1974_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1889_load_0 ptr_deref_1922_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1889_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1922_load_0_req_0;
      ptr_deref_1889_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1922_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1889_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1922_load_0_req_1;
      ptr_deref_1889_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1922_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1889_word_address_0 & ptr_deref_1922_word_address_0;
      ptr_deref_1889_data_0 <= data_out(31 downto 16);
      ptr_deref_1922_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1905_load_0 ptr_deref_1938_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1905_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1938_load_0_req_0;
      ptr_deref_1905_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1938_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1905_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1938_load_0_req_1;
      ptr_deref_1905_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1938_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1905_word_address_0 & ptr_deref_1938_word_address_0;
      ptr_deref_1905_data_0 <= data_out(63 downto 32);
      ptr_deref_1938_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1950_load_0 ptr_deref_1962_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1950_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1962_load_0_req_0;
      ptr_deref_1950_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1962_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1950_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1962_load_0_req_1;
      ptr_deref_1950_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1962_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1950_word_address_0 & ptr_deref_1962_word_address_0;
      ptr_deref_1950_data_0 <= data_out(63 downto 32);
      ptr_deref_1962_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2169_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2169_load_0_req_0;
      ptr_deref_2169_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2169_load_0_req_1;
      ptr_deref_2169_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2169_word_address_0;
      ptr_deref_2169_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2199_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2199_store_0_req_0;
      ptr_deref_2199_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2199_store_0_req_1;
      ptr_deref_2199_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2199_word_address_0;
      data_in <= ptr_deref_2199_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1844_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_start_1844_inst_req_0;
      RPIPE_Block1_start_1844_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_start_1844_inst_req_1;
      RPIPE_Block1_start_1844_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1845 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2305_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2305_inst_req_0;
      WPIPE_Block1_done_2305_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2305_inst_req_1;
      WPIPE_Block1_done_2305_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1845;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_6620_start: Boolean;
  signal convTransposeC_CP_6620_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2472_inst_req_1 : boolean;
  signal addr_of_2667_final_reg_req_1 : boolean;
  signal ptr_deref_2421_load_0_req_1 : boolean;
  signal type_cast_2472_inst_ack_1 : boolean;
  signal addr_of_2667_final_reg_ack_0 : boolean;
  signal type_cast_2472_inst_req_0 : boolean;
  signal type_cast_2599_inst_req_1 : boolean;
  signal type_cast_2472_inst_ack_0 : boolean;
  signal addr_of_2636_final_reg_req_1 : boolean;
  signal addr_of_2636_final_reg_ack_0 : boolean;
  signal ptr_deref_2445_load_0_ack_0 : boolean;
  signal addr_of_2636_final_reg_req_0 : boolean;
  signal type_cast_2599_inst_ack_1 : boolean;
  signal ptr_deref_2640_load_0_req_0 : boolean;
  signal ptr_deref_2640_load_0_ack_0 : boolean;
  signal array_obj_ref_2666_index_offset_req_0 : boolean;
  signal type_cast_2477_inst_ack_1 : boolean;
  signal type_cast_2676_inst_ack_1 : boolean;
  signal type_cast_2676_inst_req_1 : boolean;
  signal if_stmt_2689_branch_ack_1 : boolean;
  signal ptr_deref_2421_load_0_ack_1 : boolean;
  signal addr_of_2636_final_reg_ack_1 : boolean;
  signal type_cast_2676_inst_req_0 : boolean;
  signal type_cast_2676_inst_ack_0 : boolean;
  signal array_obj_ref_2635_index_offset_req_0 : boolean;
  signal array_obj_ref_2635_index_offset_ack_0 : boolean;
  signal ptr_deref_2670_store_0_req_1 : boolean;
  signal ptr_deref_2670_store_0_ack_1 : boolean;
  signal type_cast_2629_inst_req_0 : boolean;
  signal type_cast_2629_inst_ack_0 : boolean;
  signal array_obj_ref_2635_index_offset_req_1 : boolean;
  signal array_obj_ref_2666_index_offset_req_1 : boolean;
  signal array_obj_ref_2666_index_offset_ack_1 : boolean;
  signal ptr_deref_2640_load_0_req_1 : boolean;
  signal ptr_deref_2640_load_0_ack_1 : boolean;
  signal ptr_deref_2433_load_0_req_1 : boolean;
  signal type_cast_2660_inst_req_0 : boolean;
  signal if_stmt_2689_branch_req_0 : boolean;
  signal array_obj_ref_2635_index_offset_ack_1 : boolean;
  signal type_cast_2477_inst_req_0 : boolean;
  signal type_cast_2477_inst_ack_0 : boolean;
  signal ptr_deref_2670_store_0_req_0 : boolean;
  signal ptr_deref_2670_store_0_ack_0 : boolean;
  signal ptr_deref_2445_load_0_req_1 : boolean;
  signal ptr_deref_2433_load_0_ack_1 : boolean;
  signal type_cast_2660_inst_ack_0 : boolean;
  signal ptr_deref_2445_load_0_ack_1 : boolean;
  signal addr_of_2667_final_reg_req_0 : boolean;
  signal type_cast_2629_inst_req_1 : boolean;
  signal array_obj_ref_2666_index_offset_ack_0 : boolean;
  signal addr_of_2667_final_reg_ack_1 : boolean;
  signal type_cast_2629_inst_ack_1 : boolean;
  signal ptr_deref_2445_load_0_req_0 : boolean;
  signal type_cast_2660_inst_ack_1 : boolean;
  signal type_cast_2660_inst_req_1 : boolean;
  signal if_stmt_2689_branch_ack_0 : boolean;
  signal ptr_deref_2421_load_0_req_0 : boolean;
  signal type_cast_2599_inst_ack_0 : boolean;
  signal type_cast_2599_inst_req_0 : boolean;
  signal type_cast_2477_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2315_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2315_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2315_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2315_inst_ack_1 : boolean;
  signal ptr_deref_2328_load_0_req_0 : boolean;
  signal ptr_deref_2328_load_0_ack_0 : boolean;
  signal ptr_deref_2328_load_0_req_1 : boolean;
  signal ptr_deref_2328_load_0_ack_1 : boolean;
  signal type_cast_2338_inst_req_0 : boolean;
  signal type_cast_2338_inst_ack_0 : boolean;
  signal type_cast_2338_inst_req_1 : boolean;
  signal type_cast_2338_inst_ack_1 : boolean;
  signal ptr_deref_2350_load_0_req_0 : boolean;
  signal ptr_deref_2350_load_0_ack_0 : boolean;
  signal ptr_deref_2350_load_0_req_1 : boolean;
  signal ptr_deref_2350_load_0_ack_1 : boolean;
  signal ptr_deref_2362_load_0_req_0 : boolean;
  signal ptr_deref_2362_load_0_ack_0 : boolean;
  signal ptr_deref_2362_load_0_req_1 : boolean;
  signal ptr_deref_2362_load_0_ack_1 : boolean;
  signal ptr_deref_2372_load_0_req_0 : boolean;
  signal ptr_deref_2372_load_0_ack_0 : boolean;
  signal ptr_deref_2372_load_0_req_1 : boolean;
  signal ptr_deref_2372_load_0_ack_1 : boolean;
  signal type_cast_2376_inst_req_0 : boolean;
  signal type_cast_2376_inst_ack_0 : boolean;
  signal type_cast_2376_inst_req_1 : boolean;
  signal type_cast_2376_inst_ack_1 : boolean;
  signal ptr_deref_2433_load_0_ack_0 : boolean;
  signal ptr_deref_2388_load_0_req_0 : boolean;
  signal ptr_deref_2388_load_0_ack_0 : boolean;
  signal ptr_deref_2421_load_0_ack_0 : boolean;
  signal ptr_deref_2433_load_0_req_0 : boolean;
  signal ptr_deref_2388_load_0_req_1 : boolean;
  signal ptr_deref_2388_load_0_ack_1 : boolean;
  signal LOAD_padding_2391_load_0_req_0 : boolean;
  signal LOAD_padding_2391_load_0_ack_0 : boolean;
  signal LOAD_padding_2391_load_0_req_1 : boolean;
  signal LOAD_padding_2391_load_0_ack_1 : boolean;
  signal type_cast_2395_inst_req_0 : boolean;
  signal type_cast_2395_inst_ack_0 : boolean;
  signal type_cast_2395_inst_req_1 : boolean;
  signal type_cast_2395_inst_ack_1 : boolean;
  signal ptr_deref_2405_load_0_req_0 : boolean;
  signal ptr_deref_2405_load_0_ack_0 : boolean;
  signal ptr_deref_2405_load_0_req_1 : boolean;
  signal ptr_deref_2405_load_0_ack_1 : boolean;
  signal type_cast_2409_inst_req_0 : boolean;
  signal type_cast_2409_inst_ack_0 : boolean;
  signal type_cast_2409_inst_req_1 : boolean;
  signal type_cast_2409_inst_ack_1 : boolean;
  signal type_cast_2713_inst_req_0 : boolean;
  signal type_cast_2713_inst_ack_0 : boolean;
  signal type_cast_2713_inst_req_1 : boolean;
  signal type_cast_2713_inst_ack_1 : boolean;
  signal type_cast_2722_inst_req_0 : boolean;
  signal type_cast_2722_inst_ack_0 : boolean;
  signal type_cast_2722_inst_req_1 : boolean;
  signal type_cast_2722_inst_ack_1 : boolean;
  signal type_cast_2739_inst_req_0 : boolean;
  signal type_cast_2739_inst_ack_0 : boolean;
  signal type_cast_2739_inst_req_1 : boolean;
  signal type_cast_2739_inst_ack_1 : boolean;
  signal if_stmt_2746_branch_req_0 : boolean;
  signal if_stmt_2746_branch_ack_1 : boolean;
  signal if_stmt_2746_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2754_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2754_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2754_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2754_inst_ack_1 : boolean;
  signal phi_stmt_2455_req_0 : boolean;
  signal type_cast_2465_inst_req_0 : boolean;
  signal type_cast_2465_inst_ack_0 : boolean;
  signal type_cast_2465_inst_req_1 : boolean;
  signal type_cast_2465_inst_ack_1 : boolean;
  signal phi_stmt_2462_req_0 : boolean;
  signal type_cast_2461_inst_req_0 : boolean;
  signal type_cast_2461_inst_ack_0 : boolean;
  signal type_cast_2461_inst_req_1 : boolean;
  signal type_cast_2461_inst_ack_1 : boolean;
  signal phi_stmt_2455_req_1 : boolean;
  signal type_cast_2467_inst_req_0 : boolean;
  signal type_cast_2467_inst_ack_0 : boolean;
  signal type_cast_2467_inst_req_1 : boolean;
  signal type_cast_2467_inst_ack_1 : boolean;
  signal phi_stmt_2462_req_1 : boolean;
  signal phi_stmt_2455_ack_0 : boolean;
  signal phi_stmt_2462_ack_0 : boolean;
  signal type_cast_2589_inst_req_0 : boolean;
  signal type_cast_2589_inst_ack_0 : boolean;
  signal type_cast_2589_inst_req_1 : boolean;
  signal type_cast_2589_inst_ack_1 : boolean;
  signal phi_stmt_2583_req_1 : boolean;
  signal phi_stmt_2583_req_0 : boolean;
  signal phi_stmt_2583_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_6620_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6620_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_6620_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6620_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_6620: Block -- control-path 
    signal convTransposeC_CP_6620_elements: BooleanArray(92 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_6620_elements(0) <= convTransposeC_CP_6620_start;
    convTransposeC_CP_6620_symbol <= convTransposeC_CP_6620_elements(70);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2313/$entry
      -- CP-element group 0: 	 branch_block_stmt_2313/branch_block_stmt_2313__entry__
      -- CP-element group 0: 	 branch_block_stmt_2313/assign_stmt_2316__entry__
      -- CP-element group 0: 	 branch_block_stmt_2313/assign_stmt_2316/$entry
      -- CP-element group 0: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_Sample/rr
      -- 
    rr_6668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(0), ack => RPIPE_Block2_start_2315_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_Update/cr
      -- 
    ra_6669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2315_inst_ack_0, ack => convTransposeC_CP_6620_elements(1)); -- 
    cr_6673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(1), ack => RPIPE_Block2_start_2315_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2316__exit__
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452__entry__
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2316/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2316/RPIPE_Block2_start_2315_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Sample/word_access_start/$entry
      -- 
    ca_6674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2315_inst_ack_1, ack => convTransposeC_CP_6620_elements(2)); -- 
    cr_7110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2421_load_0_req_1); -- 
    cr_7160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2433_load_0_req_1); -- 
    cr_7210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2445_load_0_req_1); -- 
    rr_7199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2445_load_0_req_0); -- 
    rr_7099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2421_load_0_req_0); -- 
    rr_6710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2328_load_0_req_0); -- 
    cr_6721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2328_load_0_req_1); -- 
    cr_6740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => type_cast_2338_inst_req_1); -- 
    rr_6774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2350_load_0_req_0); -- 
    cr_6785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2350_load_0_req_1); -- 
    rr_6824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2362_load_0_req_0); -- 
    cr_6835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2362_load_0_req_1); -- 
    rr_6874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2372_load_0_req_0); -- 
    cr_6885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2372_load_0_req_1); -- 
    cr_6904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => type_cast_2376_inst_req_1); -- 
    rr_6938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2388_load_0_req_0); -- 
    rr_7149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2433_load_0_req_0); -- 
    cr_6949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2388_load_0_req_1); -- 
    rr_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => LOAD_padding_2391_load_0_req_0); -- 
    cr_6982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => LOAD_padding_2391_load_0_req_1); -- 
    cr_7001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => type_cast_2395_inst_req_1); -- 
    rr_7035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2405_load_0_req_0); -- 
    cr_7046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => ptr_deref_2405_load_0_req_1); -- 
    cr_7065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(2), ack => type_cast_2409_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Sample/word_access_start/word_0/ra
      -- 
    ra_6711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2328_load_0_ack_0, ack => convTransposeC_CP_6620_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/ptr_deref_2328_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/ptr_deref_2328_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/ptr_deref_2328_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2328_Update/ptr_deref_2328_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_Sample/rr
      -- 
    ca_6722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2328_load_0_ack_1, ack => convTransposeC_CP_6620_elements(4)); -- 
    rr_6735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(4), ack => type_cast_2338_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_Sample/ra
      -- 
    ra_6736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2338_inst_ack_0, ack => convTransposeC_CP_6620_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2338_Update/ca
      -- 
    ca_6741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2338_inst_ack_1, ack => convTransposeC_CP_6620_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Sample/word_access_start/word_0/ra
      -- 
    ra_6775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2350_load_0_ack_0, ack => convTransposeC_CP_6620_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/ptr_deref_2350_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/ptr_deref_2350_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/ptr_deref_2350_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2350_Update/ptr_deref_2350_Merge/merge_ack
      -- 
    ca_6786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2350_load_0_ack_1, ack => convTransposeC_CP_6620_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Sample/word_access_start/word_0/ra
      -- 
    ra_6825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2362_load_0_ack_0, ack => convTransposeC_CP_6620_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	31 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/ptr_deref_2362_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/ptr_deref_2362_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/ptr_deref_2362_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2362_Update/ptr_deref_2362_Merge/merge_ack
      -- 
    ca_6836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2362_load_0_ack_1, ack => convTransposeC_CP_6620_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Sample/word_access_start/word_0/ra
      -- 
    ra_6875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2372_load_0_ack_0, ack => convTransposeC_CP_6620_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (12) 
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/ptr_deref_2372_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/ptr_deref_2372_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/ptr_deref_2372_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2372_Update/ptr_deref_2372_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_Sample/rr
      -- 
    ca_6886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2372_load_0_ack_1, ack => convTransposeC_CP_6620_elements(12)); -- 
    rr_6899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(12), ack => type_cast_2376_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_Sample/ra
      -- 
    ra_6900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2376_inst_ack_0, ack => convTransposeC_CP_6620_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2376_Update/ca
      -- 
    ca_6905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2376_inst_ack_1, ack => convTransposeC_CP_6620_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Sample/word_access_start/word_0/ra
      -- 
    ra_6939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2388_load_0_ack_0, ack => convTransposeC_CP_6620_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/ptr_deref_2388_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/ptr_deref_2388_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/ptr_deref_2388_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2388_Update/ptr_deref_2388_Merge/merge_ack
      -- 
    ca_6950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2388_load_0_ack_1, ack => convTransposeC_CP_6620_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Sample/word_access_start/word_0/ra
      -- 
    ra_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2391_load_0_ack_0, ack => convTransposeC_CP_6620_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/LOAD_padding_2391_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/LOAD_padding_2391_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/LOAD_padding_2391_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/LOAD_padding_2391_Update/LOAD_padding_2391_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_Sample/rr
      -- 
    ca_6983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2391_load_0_ack_1, ack => convTransposeC_CP_6620_elements(18)); -- 
    rr_6996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(18), ack => type_cast_2395_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_Sample/ra
      -- 
    ra_6997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2395_inst_ack_0, ack => convTransposeC_CP_6620_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	31 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2395_Update/ca
      -- 
    ca_7002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2395_inst_ack_1, ack => convTransposeC_CP_6620_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Sample/word_access_start/word_0/ra
      -- 
    ra_7036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2405_load_0_ack_0, ack => convTransposeC_CP_6620_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (12) 
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/ptr_deref_2405_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/ptr_deref_2405_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/ptr_deref_2405_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2405_Update/ptr_deref_2405_Merge/merge_ack
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_Sample/rr
      -- 
    ca_7047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2405_load_0_ack_1, ack => convTransposeC_CP_6620_elements(22)); -- 
    rr_7060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(22), ack => type_cast_2409_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_Sample/ra
      -- 
    ra_7061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2409_inst_ack_0, ack => convTransposeC_CP_6620_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/type_cast_2409_Update/ca
      -- 
    ca_7066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2409_inst_ack_1, ack => convTransposeC_CP_6620_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Sample/word_access_start/$exit
      -- 
    ra_7100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2421_load_0_ack_0, ack => convTransposeC_CP_6620_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/ptr_deref_2421_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/ptr_deref_2421_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/ptr_deref_2421_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_Update/ptr_deref_2421_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2421_update_completed_
      -- 
    ca_7111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2421_load_0_ack_1, ack => convTransposeC_CP_6620_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Sample/word_access_start/word_0/ra
      -- 
    ra_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2433_load_0_ack_0, ack => convTransposeC_CP_6620_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/ptr_deref_2433_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/ptr_deref_2433_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/ptr_deref_2433_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2433_Update/ptr_deref_2433_Merge/merge_ack
      -- 
    ca_7161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2433_load_0_ack_1, ack => convTransposeC_CP_6620_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Sample/word_access_start/word_0/ra
      -- CP-element group 29: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_sample_completed_
      -- 
    ra_7200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2445_load_0_ack_0, ack => convTransposeC_CP_6620_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/ptr_deref_2445_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/ptr_deref_2445_Merge/merge_ack
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/ptr_deref_2445_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/ptr_deref_2445_Update/ptr_deref_2445_Merge/$exit
      -- 
    ca_7211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2445_load_0_ack_1, ack => convTransposeC_CP_6620_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	10 
    -- CP-element group 31: 	20 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	6 
    -- CP-element group 31: 	8 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	71 
    -- CP-element group 31: 	72 
    -- CP-element group 31: 	73 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452/$exit
      -- CP-element group 31: 	 branch_block_stmt_2313/assign_stmt_2325_to_assign_stmt_2452__exit__
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/Update/cr
      -- 
    rr_7628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(31), ack => type_cast_2465_inst_req_0); -- 
    cr_7633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(31), ack => type_cast_2465_inst_req_1); -- 
    convTransposeC_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(10) & convTransposeC_CP_6620_elements(20) & convTransposeC_CP_6620_elements(26) & convTransposeC_CP_6620_elements(30) & convTransposeC_CP_6620_elements(14) & convTransposeC_CP_6620_elements(24) & convTransposeC_CP_6620_elements(28) & convTransposeC_CP_6620_elements(16) & convTransposeC_CP_6620_elements(6) & convTransposeC_CP_6620_elements(8);
      gj_convTransposeC_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	86 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_sample_completed_
      -- 
    ra_7228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2472_inst_ack_0, ack => convTransposeC_CP_6620_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	86 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_update_completed_
      -- 
    ca_7233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2472_inst_ack_1, ack => convTransposeC_CP_6620_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	86 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_Sample/ra
      -- 
    ra_7242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2477_inst_ack_0, ack => convTransposeC_CP_6620_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	86 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_Update/$exit
      -- 
    ca_7247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2477_inst_ack_1, ack => convTransposeC_CP_6620_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	90 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580__exit__
      -- CP-element group 36: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/$exit
      -- CP-element group 36: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2583/$entry
      -- CP-element group 36: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/$entry
      -- 
    convTransposeC_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(33) & convTransposeC_CP_6620_elements(35);
      gj_convTransposeC_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_Sample/$exit
      -- 
    ra_7259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2599_inst_ack_0, ack => convTransposeC_CP_6620_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	92 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_Update/$exit
      -- 
    ca_7264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2599_inst_ack_1, ack => convTransposeC_CP_6620_elements(38)); -- 
    rr_7272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(38), ack => type_cast_2629_inst_req_0); -- 
    rr_7382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(38), ack => type_cast_2660_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_Sample/ra
      -- 
    ra_7273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2629_inst_ack_0, ack => convTransposeC_CP_6620_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	92 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_Sample/req
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_index_resize_1/index_resize_req
      -- 
    ca_7278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2629_inst_ack_1, ack => convTransposeC_CP_6620_elements(40)); -- 
    req_7303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(40), ack => array_obj_ref_2635_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_Sample/ack
      -- 
    ack_7304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2635_index_offset_ack_0, ack => convTransposeC_CP_6620_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	92 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_request/req
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_request/$entry
      -- 
    ack_7309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2635_index_offset_ack_1, ack => convTransposeC_CP_6620_elements(42)); -- 
    req_7318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(42), ack => addr_of_2636_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_request/ack
      -- CP-element group 43: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_sample_completed_
      -- 
    ack_7319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2636_final_reg_ack_0, ack => convTransposeC_CP_6620_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	92 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Sample/word_access_start/word_0/rr
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_base_address_calculated
      -- 
    ack_7324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2636_final_reg_ack_1, ack => convTransposeC_CP_6620_elements(44)); -- 
    rr_7357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(44), ack => ptr_deref_2640_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Sample/word_access_start/word_0/ra
      -- CP-element group 45: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_sample_completed_
      -- 
    ra_7358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_load_0_ack_0, ack => convTransposeC_CP_6620_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/ptr_deref_2640_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/ptr_deref_2640_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/ptr_deref_2640_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/ptr_deref_2640_Merge/merge_ack
      -- CP-element group 46: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_update_completed_
      -- 
    ca_7369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_load_0_ack_1, ack => convTransposeC_CP_6620_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_Sample/ra
      -- 
    ra_7383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2660_inst_ack_0, ack => convTransposeC_CP_6620_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	92 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_Sample/req
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_Update/ca
      -- 
    ca_7388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2660_inst_ack_1, ack => convTransposeC_CP_6620_elements(48)); -- 
    req_7413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(48), ack => array_obj_ref_2666_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_Sample/ack
      -- 
    ack_7414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2666_index_offset_ack_0, ack => convTransposeC_CP_6620_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	92 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_request/req
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_root_address_calculated
      -- 
    ack_7419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2666_index_offset_ack_1, ack => convTransposeC_CP_6620_elements(50)); -- 
    req_7428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(50), ack => addr_of_2667_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_request/ack
      -- CP-element group 51: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_request/$exit
      -- 
    ack_7429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2667_final_reg_ack_0, ack => convTransposeC_CP_6620_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	92 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_complete/ack
      -- 
    ack_7434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2667_final_reg_ack_1, ack => convTransposeC_CP_6620_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/ptr_deref_2670_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/ptr_deref_2670_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/ptr_deref_2670_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/ptr_deref_2670_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/word_access_start/word_0/rr
      -- CP-element group 53: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_sample_start_
      -- 
    rr_7472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(53), ack => ptr_deref_2670_store_0_req_0); -- 
    convTransposeC_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(46) & convTransposeC_CP_6620_elements(52);
      gj_convTransposeC_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/word_access_start/word_0/ra
      -- CP-element group 54: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_sample_completed_
      -- 
    ra_7473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2670_store_0_ack_0, ack => convTransposeC_CP_6620_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	92 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_update_completed_
      -- 
    ca_7484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2670_store_0_ack_1, ack => convTransposeC_CP_6620_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	92 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_Sample/$exit
      -- 
    ra_7493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2676_inst_ack_0, ack => convTransposeC_CP_6620_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	92 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_update_completed_
      -- 
    ca_7498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2676_inst_ack_1, ack => convTransposeC_CP_6620_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_2313/if_stmt_2689_else_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2313/if_stmt_2689_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/$exit
      -- CP-element group 58: 	 branch_block_stmt_2313/if_stmt_2689_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_2313/if_stmt_2689_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_2313/if_stmt_2689_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_2313/if_stmt_2689_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688__exit__
      -- CP-element group 58: 	 branch_block_stmt_2313/if_stmt_2689__entry__
      -- CP-element group 58: 	 branch_block_stmt_2313/R_cmp_2690_place
      -- 
    branch_req_7506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(58), ack => if_stmt_2689_branch_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(57) & convTransposeC_CP_6620_elements(41) & convTransposeC_CP_6620_elements(55) & convTransposeC_CP_6620_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	87 
    -- CP-element group 59: 	88 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_2313/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_2313/if_stmt_2689_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_2313/if_stmt_2689_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_2313/merge_stmt_2695__exit__
      -- CP-element group 59: 	 branch_block_stmt_2313/assign_stmt_2701__entry__
      -- CP-element group 59: 	 branch_block_stmt_2313/assign_stmt_2701__exit__
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_2313/assign_stmt_2701/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/assign_stmt_2701/$exit
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_2313/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_2313/merge_stmt_2695_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_2313/merge_stmt_2695_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_2313/merge_stmt_2695_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_2313/merge_stmt_2695_PhiAck/dummy
      -- 
    if_choice_transition_7511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2689_branch_ack_1, ack => convTransposeC_CP_6620_elements(59)); -- 
    rr_7709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(59), ack => type_cast_2589_inst_req_0); -- 
    cr_7714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(59), ack => type_cast_2589_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60: 	64 
    -- CP-element group 60: 	66 
    -- CP-element group 60:  members (24) 
      -- CP-element group 60: 	 branch_block_stmt_2313/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_2313/if_stmt_2689_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_2313/if_stmt_2689_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_2313/merge_stmt_2703__exit__
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745__entry__
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/$entry
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2313/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_2313/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_2313/merge_stmt_2703_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_2313/merge_stmt_2703_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_2313/merge_stmt_2703_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_2313/merge_stmt_2703_PhiAck/dummy
      -- 
    else_choice_transition_7515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2689_branch_ack_0, ack => convTransposeC_CP_6620_elements(60)); -- 
    rr_7531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(60), ack => type_cast_2713_inst_req_0); -- 
    cr_7536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(60), ack => type_cast_2713_inst_req_1); -- 
    cr_7550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(60), ack => type_cast_2722_inst_req_1); -- 
    cr_7564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(60), ack => type_cast_2739_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_Sample/ra
      -- 
    ra_7532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2713_inst_ack_0, ack => convTransposeC_CP_6620_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2713_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_Sample/rr
      -- 
    ca_7537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2713_inst_ack_1, ack => convTransposeC_CP_6620_elements(62)); -- 
    rr_7545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(62), ack => type_cast_2722_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_Sample/ra
      -- 
    ra_7546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_0, ack => convTransposeC_CP_6620_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	60 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2722_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_Sample/rr
      -- 
    ca_7551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_1, ack => convTransposeC_CP_6620_elements(64)); -- 
    rr_7559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(64), ack => type_cast_2739_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_Sample/ra
      -- 
    ra_7560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2739_inst_ack_0, ack => convTransposeC_CP_6620_elements(65)); -- 
    -- CP-element group 66:  branch  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (13) 
      -- CP-element group 66: 	 branch_block_stmt_2313/R_cmp87_2747_place
      -- CP-element group 66: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745__exit__
      -- CP-element group 66: 	 branch_block_stmt_2313/if_stmt_2746__entry__
      -- CP-element group 66: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/$exit
      -- CP-element group 66: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2313/assign_stmt_2709_to_assign_stmt_2745/type_cast_2739_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_2313/if_stmt_2746_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2313/if_stmt_2746_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2313/if_stmt_2746_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2313/if_stmt_2746_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2313/if_stmt_2746_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2313/if_stmt_2746_else_link/$entry
      -- 
    ca_7565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2739_inst_ack_1, ack => convTransposeC_CP_6620_elements(66)); -- 
    branch_req_7573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(66), ack => if_stmt_2746_branch_req_0); -- 
    -- CP-element group 67:  merge  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (15) 
      -- CP-element group 67: 	 branch_block_stmt_2313/ifx_xelse_whilex_xend
      -- CP-element group 67: 	 branch_block_stmt_2313/merge_stmt_2752__exit__
      -- CP-element group 67: 	 branch_block_stmt_2313/assign_stmt_2756__entry__
      -- CP-element group 67: 	 branch_block_stmt_2313/if_stmt_2746_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2313/if_stmt_2746_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2313/assign_stmt_2756/$entry
      -- CP-element group 67: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_2313/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2313/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2313/merge_stmt_2752_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2313/merge_stmt_2752_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2313/merge_stmt_2752_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2313/merge_stmt_2752_PhiAck/dummy
      -- 
    if_choice_transition_7578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2746_branch_ack_1, ack => convTransposeC_CP_6620_elements(67)); -- 
    req_7595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(67), ack => WPIPE_Block2_done_2754_inst_req_0); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	76 
    -- CP-element group 68: 	77 
    -- CP-element group 68: 	79 
    -- CP-element group 68: 	80 
    -- CP-element group 68:  members (20) 
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 68: 	 branch_block_stmt_2313/if_stmt_2746_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2313/if_stmt_2746_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2746_branch_ack_0, ack => convTransposeC_CP_6620_elements(68)); -- 
    rr_7654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(68), ack => type_cast_2461_inst_req_0); -- 
    cr_7659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(68), ack => type_cast_2461_inst_req_1); -- 
    rr_7677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(68), ack => type_cast_2467_inst_req_0); -- 
    cr_7682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(68), ack => type_cast_2467_inst_req_1); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_update_start_
      -- CP-element group 69: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_Update/req
      -- 
    ack_7596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2754_inst_ack_0, ack => convTransposeC_CP_6620_elements(69)); -- 
    req_7600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(69), ack => WPIPE_Block2_done_2754_inst_req_1); -- 
    -- CP-element group 70:  transition  place  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (16) 
      -- CP-element group 70: 	 $exit
      -- CP-element group 70: 	 branch_block_stmt_2313/$exit
      -- CP-element group 70: 	 branch_block_stmt_2313/branch_block_stmt_2313__exit__
      -- CP-element group 70: 	 branch_block_stmt_2313/assign_stmt_2756__exit__
      -- CP-element group 70: 	 branch_block_stmt_2313/return__
      -- CP-element group 70: 	 branch_block_stmt_2313/merge_stmt_2758__exit__
      -- CP-element group 70: 	 branch_block_stmt_2313/assign_stmt_2756/$exit
      -- CP-element group 70: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2313/assign_stmt_2756/WPIPE_Block2_done_2754_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_2313/return___PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2313/return___PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2313/merge_stmt_2758_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2313/merge_stmt_2758_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2313/merge_stmt_2758_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2313/merge_stmt_2758_PhiAck/dummy
      -- 
    ack_7601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2754_inst_ack_1, ack => convTransposeC_CP_6620_elements(70)); -- 
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/$exit
      -- CP-element group 71: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2459_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_req
      -- 
    phi_stmt_2455_req_7612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2455_req_7612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(71), ack => phi_stmt_2455_req_0); -- 
    -- Element group convTransposeC_CP_6620_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_6620_elements(31), ack => convTransposeC_CP_6620_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	31 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/Sample/ra
      -- 
    ra_7629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2465_inst_ack_0, ack => convTransposeC_CP_6620_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/Update/ca
      -- 
    ca_7634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2465_inst_ack_1, ack => convTransposeC_CP_6620_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/$exit
      -- CP-element group 74: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/$exit
      -- CP-element group 74: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2465/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_req
      -- 
    phi_stmt_2462_req_7635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2462_req_7635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(74), ack => phi_stmt_2462_req_0); -- 
    convTransposeC_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(72) & convTransposeC_CP_6620_elements(73);
      gj_convTransposeC_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	83 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2313/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(71) & convTransposeC_CP_6620_elements(74);
      gj_convTransposeC_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	68 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Sample/ra
      -- 
    ra_7655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2461_inst_ack_0, ack => convTransposeC_CP_6620_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	68 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/Update/ca
      -- 
    ca_7660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2461_inst_ack_1, ack => convTransposeC_CP_6620_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	82 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/$exit
      -- CP-element group 78: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/$exit
      -- CP-element group 78: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2461/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2455/phi_stmt_2455_req
      -- 
    phi_stmt_2455_req_7661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2455_req_7661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(78), ack => phi_stmt_2455_req_1); -- 
    convTransposeC_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(76) & convTransposeC_CP_6620_elements(77);
      gj_convTransposeC_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	68 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/Sample/ra
      -- 
    ra_7678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2467_inst_ack_0, ack => convTransposeC_CP_6620_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	68 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/Update/ca
      -- 
    ca_7683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2467_inst_ack_1, ack => convTransposeC_CP_6620_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/$exit
      -- CP-element group 81: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/$exit
      -- CP-element group 81: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_sources/type_cast_2467/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2462/phi_stmt_2462_req
      -- 
    phi_stmt_2462_req_7684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2462_req_7684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(81), ack => phi_stmt_2462_req_1); -- 
    convTransposeC_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(79) & convTransposeC_CP_6620_elements(80);
      gj_convTransposeC_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2313/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(78) & convTransposeC_CP_6620_elements(81);
      gj_convTransposeC_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  merge  fork  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	75 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2313/merge_stmt_2454_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_2313/merge_stmt_2454_PhiAck/$entry
      -- 
    convTransposeC_CP_6620_elements(83) <= OrReduce(convTransposeC_CP_6620_elements(75) & convTransposeC_CP_6620_elements(82));
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2313/merge_stmt_2454_PhiAck/phi_stmt_2455_ack
      -- 
    phi_stmt_2455_ack_7689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2455_ack_0, ack => convTransposeC_CP_6620_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2313/merge_stmt_2454_PhiAck/phi_stmt_2462_ack
      -- 
    phi_stmt_2462_ack_7690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2462_ack_0, ack => convTransposeC_CP_6620_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	32 
    -- CP-element group 86: 	33 
    -- CP-element group 86: 	34 
    -- CP-element group 86: 	35 
    -- CP-element group 86:  members (16) 
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2472_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/type_cast_2477_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2313/merge_stmt_2454__exit__
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580__entry__
      -- CP-element group 86: 	 branch_block_stmt_2313/assign_stmt_2473_to_assign_stmt_2580/$entry
      -- CP-element group 86: 	 branch_block_stmt_2313/merge_stmt_2454_PhiAck/$exit
      -- 
    cr_7232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(86), ack => type_cast_2472_inst_req_1); -- 
    rr_7227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(86), ack => type_cast_2472_inst_req_0); -- 
    rr_7241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(86), ack => type_cast_2477_inst_req_0); -- 
    cr_7246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(86), ack => type_cast_2477_inst_req_1); -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(84) & convTransposeC_CP_6620_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	59 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/Sample/ra
      -- 
    ra_7710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_0, ack => convTransposeC_CP_6620_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	59 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/Update/ca
      -- 
    ca_7715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_1, ack => convTransposeC_CP_6620_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/$exit
      -- CP-element group 89: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/$exit
      -- CP-element group 89: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2589/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_2313/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_req
      -- 
    phi_stmt_2583_req_7716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2583_req_7716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(89), ack => phi_stmt_2583_req_1); -- 
    convTransposeC_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6620_elements(87) & convTransposeC_CP_6620_elements(88);
      gj_convTransposeC_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6620_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  output  delay-element  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	36 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2583/$exit
      -- CP-element group 90: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_sources/type_cast_2587_konst_delay_trans
      -- CP-element group 90: 	 branch_block_stmt_2313/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2583/phi_stmt_2583_req
      -- 
    phi_stmt_2583_req_7727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2583_req_7727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(90), ack => phi_stmt_2583_req_0); -- 
    -- Element group convTransposeC_CP_6620_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => convTransposeC_CP_6620_elements(36), ack => convTransposeC_CP_6620_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  merge  transition  place  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2313/merge_stmt_2582_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_2313/merge_stmt_2582_PhiAck/$entry
      -- 
    convTransposeC_CP_6620_elements(91) <= OrReduce(convTransposeC_CP_6620_elements(89) & convTransposeC_CP_6620_elements(90));
    -- CP-element group 92:  fork  transition  place  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	56 
    -- CP-element group 92: 	57 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	38 
    -- CP-element group 92: 	40 
    -- CP-element group 92: 	42 
    -- CP-element group 92: 	48 
    -- CP-element group 92: 	55 
    -- CP-element group 92: 	50 
    -- CP-element group 92: 	52 
    -- CP-element group 92: 	44 
    -- CP-element group 92:  members (45) 
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2636_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2676_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2635_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/array_obj_ref_2666_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/addr_of_2667_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2640_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2629_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/ptr_deref_2670_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2660_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688/type_cast_2599_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2313/merge_stmt_2582__exit__
      -- CP-element group 92: 	 branch_block_stmt_2313/assign_stmt_2596_to_assign_stmt_2688__entry__
      -- CP-element group 92: 	 branch_block_stmt_2313/merge_stmt_2582_PhiAck/$exit
      -- CP-element group 92: 	 branch_block_stmt_2313/merge_stmt_2582_PhiAck/phi_stmt_2583_ack
      -- 
    phi_stmt_2583_ack_7732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2583_ack_0, ack => convTransposeC_CP_6620_elements(92)); -- 
    req_7433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => addr_of_2667_final_reg_req_1); -- 
    cr_7263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => type_cast_2599_inst_req_1); -- 
    req_7323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => addr_of_2636_final_reg_req_1); -- 
    cr_7497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => type_cast_2676_inst_req_1); -- 
    rr_7492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => type_cast_2676_inst_req_0); -- 
    cr_7483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => ptr_deref_2670_store_0_req_1); -- 
    req_7308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => array_obj_ref_2635_index_offset_req_1); -- 
    req_7418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => array_obj_ref_2666_index_offset_req_1); -- 
    cr_7368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => ptr_deref_2640_load_0_req_1); -- 
    cr_7277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => type_cast_2629_inst_req_1); -- 
    cr_7387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => type_cast_2660_inst_req_1); -- 
    rr_7258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6620_elements(92), ack => type_cast_2599_inst_req_0); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2542_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2563_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2623_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2654_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2391_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2391_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom62_2665_resized : std_logic_vector(13 downto 0);
    signal R_idxprom62_2665_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2634_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2634_scaled : std_logic_vector(13 downto 0);
    signal add18_2605 : std_logic_vector(31 downto 0);
    signal add26_2503 : std_logic_vector(31 downto 0);
    signal add37_2518 : std_logic_vector(31 downto 0);
    signal add52_2575 : std_logic_vector(31 downto 0);
    signal add54_2610 : std_logic_vector(31 downto 0);
    signal add67_2683 : std_logic_vector(31 downto 0);
    signal add_2488 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2635_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2635_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2635_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2635_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2635_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2635_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2666_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2666_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2666_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2666_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2666_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2666_root_address : std_logic_vector(13 downto 0);
    signal arrayidx63_2668 : std_logic_vector(31 downto 0);
    signal arrayidx_2637 : std_logic_vector(31 downto 0);
    signal call_2316 : std_logic_vector(15 downto 0);
    signal cmp79_2719 : std_logic_vector(0 downto 0);
    signal cmp87_2745 : std_logic_vector(0 downto 0);
    signal cmp_2688 : std_logic_vector(0 downto 0);
    signal conv10100_2600 : std_logic_vector(31 downto 0);
    signal conv13_2473 : std_logic_vector(31 downto 0);
    signal conv16_2478 : std_logic_vector(31 downto 0);
    signal conv23_2377 : std_logic_vector(31 downto 0);
    signal conv28_2396 : std_logic_vector(31 downto 0);
    signal conv34_2410 : std_logic_vector(31 downto 0);
    signal conv47_2544 : std_logic_vector(31 downto 0);
    signal conv50_2565 : std_logic_vector(31 downto 0);
    signal conv66_2677 : std_logic_vector(31 downto 0);
    signal conv76_2714 : std_logic_vector(31 downto 0);
    signal conv85_2740 : std_logic_vector(31 downto 0);
    signal conv_2339 : std_logic_vector(15 downto 0);
    signal div78_2452 : std_logic_vector(31 downto 0);
    signal div_2335 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2442 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2325 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2347 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2359 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2369 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2385 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2402 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2418 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2430 : std_logic_vector(31 downto 0);
    signal idxprom62_2661 : std_logic_vector(63 downto 0);
    signal idxprom_2630 : std_logic_vector(63 downto 0);
    signal inc83_2723 : std_logic_vector(15 downto 0);
    signal inc83x_xinput_dim0x_x2_2728 : std_logic_vector(15 downto 0);
    signal inc_2709 : std_logic_vector(15 downto 0);
    signal indvar_2583 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2701 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2462 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2455 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2735 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2596 : std_logic_vector(15 downto 0);
    signal mul17_2493 : std_logic_vector(31 downto 0);
    signal mul24_2498 : std_logic_vector(31 downto 0);
    signal mul35_2513 : std_logic_vector(31 downto 0);
    signal mul51_2570 : std_logic_vector(31 downto 0);
    signal mul53_2580 : std_logic_vector(31 downto 0);
    signal mul_2483 : std_logic_vector(31 downto 0);
    signal ptr_deref_2328_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2328_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2328_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2328_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2328_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2350_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2350_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2350_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2350_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2350_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2362_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2362_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2362_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2362_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2362_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2372_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2372_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2372_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2372_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2372_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2388_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2388_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2388_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2388_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2388_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2405_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2405_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2405_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2405_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2405_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2421_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2421_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2421_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2421_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2421_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2433_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2433_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2433_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2433_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2433_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2445_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2445_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2445_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2445_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2445_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2640_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2640_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2640_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2640_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2640_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2670_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2670_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2670_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2670_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2670_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2670_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext101_2556 : std_logic_vector(31 downto 0);
    signal sext103_2616 : std_logic_vector(31 downto 0);
    signal sext104_2647 : std_logic_vector(31 downto 0);
    signal sext_2535 : std_logic_vector(31 downto 0);
    signal shr61_2656 : std_logic_vector(31 downto 0);
    signal shr_2625 : std_logic_vector(31 downto 0);
    signal sub29_2550 : std_logic_vector(31 downto 0);
    signal sub40_2523 : std_logic_vector(31 downto 0);
    signal sub41_2529 : std_logic_vector(31 downto 0);
    signal sub_2508 : std_logic_vector(31 downto 0);
    signal tmp11_2351 : std_logic_vector(31 downto 0);
    signal tmp14_2363 : std_logic_vector(31 downto 0);
    signal tmp22_2373 : std_logic_vector(15 downto 0);
    signal tmp25_2389 : std_logic_vector(31 downto 0);
    signal tmp27_2392 : std_logic_vector(15 downto 0);
    signal tmp33_2406 : std_logic_vector(15 downto 0);
    signal tmp36_2422 : std_logic_vector(31 downto 0);
    signal tmp45_2434 : std_logic_vector(31 downto 0);
    signal tmp48_2446 : std_logic_vector(31 downto 0);
    signal tmp58_2641 : std_logic_vector(63 downto 0);
    signal tmp_2329 : std_logic_vector(31 downto 0);
    signal type_cast_2333_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2450_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2459_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2461_wire : std_logic_vector(15 downto 0);
    signal type_cast_2465_wire : std_logic_vector(15 downto 0);
    signal type_cast_2467_wire : std_logic_vector(15 downto 0);
    signal type_cast_2471_wire : std_logic_vector(31 downto 0);
    signal type_cast_2476_wire : std_logic_vector(31 downto 0);
    signal type_cast_2527_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2533_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2538_wire : std_logic_vector(31 downto 0);
    signal type_cast_2541_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2548_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2554_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2559_wire : std_logic_vector(31 downto 0);
    signal type_cast_2562_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2587_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2589_wire : std_logic_vector(15 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2614_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2619_wire : std_logic_vector(31 downto 0);
    signal type_cast_2622_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2628_wire : std_logic_vector(63 downto 0);
    signal type_cast_2645_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2650_wire : std_logic_vector(31 downto 0);
    signal type_cast_2653_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2659_wire : std_logic_vector(63 downto 0);
    signal type_cast_2675_wire : std_logic_vector(31 downto 0);
    signal type_cast_2681_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2699_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2707_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2712_wire : std_logic_vector(31 downto 0);
    signal type_cast_2732_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2738_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2391_word_address_0 <= "0";
    array_obj_ref_2635_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2635_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2635_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2635_resized_base_address <= "00000000000000";
    array_obj_ref_2666_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2666_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2666_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2666_resized_base_address <= "00000000000000";
    iNsTr_10_2442 <= "00000000000000000000000000000011";
    iNsTr_2_2325 <= "00000000000000000000000000000010";
    iNsTr_3_2347 <= "00000000000000000000000000000100";
    iNsTr_4_2359 <= "00000000000000000000000000000011";
    iNsTr_5_2369 <= "00000000000000000000000000000000";
    iNsTr_6_2385 <= "00000000000000000000000000000011";
    iNsTr_7_2402 <= "00000000000000000000000000000001";
    iNsTr_8_2418 <= "00000000000000000000000000000100";
    iNsTr_9_2430 <= "00000000000000000000000000000100";
    ptr_deref_2328_word_offset_0 <= "0000000";
    ptr_deref_2350_word_offset_0 <= "0000000";
    ptr_deref_2362_word_offset_0 <= "0000000";
    ptr_deref_2372_word_offset_0 <= "0";
    ptr_deref_2388_word_offset_0 <= "0000000";
    ptr_deref_2405_word_offset_0 <= "0";
    ptr_deref_2421_word_offset_0 <= "0000000";
    ptr_deref_2433_word_offset_0 <= "0000000";
    ptr_deref_2445_word_offset_0 <= "0000000";
    ptr_deref_2640_word_offset_0 <= "00000000000000";
    ptr_deref_2670_word_offset_0 <= "00000000000000";
    type_cast_2333_wire_constant <= "00000000000000000000000000000001";
    type_cast_2450_wire_constant <= "00000000000000000000000000000001";
    type_cast_2459_wire_constant <= "0000000000000000";
    type_cast_2527_wire_constant <= "00000000000000000000000000010000";
    type_cast_2533_wire_constant <= "11111111111111110000000000000000";
    type_cast_2541_wire_constant <= "00000000000000000000000000010000";
    type_cast_2548_wire_constant <= "00000000000000000000000000010000";
    type_cast_2554_wire_constant <= "11111111111111110000000000000000";
    type_cast_2562_wire_constant <= "00000000000000000000000000010000";
    type_cast_2587_wire_constant <= "0000000000000000";
    type_cast_2594_wire_constant <= "0000000000000100";
    type_cast_2614_wire_constant <= "00000000000000000000000000010000";
    type_cast_2622_wire_constant <= "00000000000000000000000000010010";
    type_cast_2645_wire_constant <= "00000000000000000000000000010000";
    type_cast_2653_wire_constant <= "00000000000000000000000000010010";
    type_cast_2681_wire_constant <= "00000000000000000000000000000100";
    type_cast_2699_wire_constant <= "0000000000000001";
    type_cast_2707_wire_constant <= "0000000000000001";
    type_cast_2732_wire_constant <= "0000000000000000";
    phi_stmt_2455: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2459_wire_constant & type_cast_2461_wire;
      req <= phi_stmt_2455_req_0 & phi_stmt_2455_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2455",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2455_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2455,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2455
    phi_stmt_2462: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2465_wire & type_cast_2467_wire;
      req <= phi_stmt_2462_req_0 & phi_stmt_2462_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2462",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2462_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2462,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2462
    phi_stmt_2583: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2587_wire_constant & type_cast_2589_wire;
      req <= phi_stmt_2583_req_0 & phi_stmt_2583_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2583",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2583_ack_0,
          idata => idata,
          odata => indvar_2583,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2583
    -- flow-through select operator MUX_2734_inst
    input_dim1x_x2_2735 <= type_cast_2732_wire_constant when (cmp79_2719(0) /=  '0') else inc_2709;
    addr_of_2636_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2636_final_reg_req_0;
      addr_of_2636_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2636_final_reg_req_1;
      addr_of_2636_final_reg_ack_1<= rack(0);
      addr_of_2636_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2636_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2635_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2637,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2667_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2667_final_reg_req_0;
      addr_of_2667_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2667_final_reg_req_1;
      addr_of_2667_final_reg_ack_1<= rack(0);
      addr_of_2667_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2667_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2666_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx63_2668,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2338_inst_req_0;
      type_cast_2338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2338_inst_req_1;
      type_cast_2338_inst_ack_1<= rack(0);
      type_cast_2338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2376_inst_req_0;
      type_cast_2376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2376_inst_req_1;
      type_cast_2376_inst_ack_1<= rack(0);
      type_cast_2376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp22_2373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_2377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2395_inst_req_0;
      type_cast_2395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2395_inst_req_1;
      type_cast_2395_inst_ack_1<= rack(0);
      type_cast_2395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp27_2392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_2396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2409_inst_req_0;
      type_cast_2409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2409_inst_req_1;
      type_cast_2409_inst_ack_1<= rack(0);
      type_cast_2409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp33_2406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_2410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2461_inst_req_0;
      type_cast_2461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2461_inst_req_1;
      type_cast_2461_inst_ack_1<= rack(0);
      type_cast_2461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2461_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2465_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2465_inst_req_0;
      type_cast_2465_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2465_inst_req_1;
      type_cast_2465_inst_ack_1<= rack(0);
      type_cast_2465_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2465_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2465_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2467_inst_req_0;
      type_cast_2467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2467_inst_req_1;
      type_cast_2467_inst_ack_1<= rack(0);
      type_cast_2467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc83x_xinput_dim0x_x2_2728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2467_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2472_inst_req_0;
      type_cast_2472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2472_inst_req_1;
      type_cast_2472_inst_ack_1<= rack(0);
      type_cast_2472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2471_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_2473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2477_inst_req_0;
      type_cast_2477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2477_inst_req_1;
      type_cast_2477_inst_ack_1<= rack(0);
      type_cast_2477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2476_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2538_inst
    process(sext_2535) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2535(31 downto 0);
      type_cast_2538_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2543_inst
    process(ASHR_i32_i32_2542_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2542_wire(31 downto 0);
      conv47_2544 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2559_inst
    process(sext101_2556) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext101_2556(31 downto 0);
      type_cast_2559_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2564_inst
    process(ASHR_i32_i32_2563_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2563_wire(31 downto 0);
      conv50_2565 <= tmp_var; -- 
    end process;
    type_cast_2589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2589_inst_req_0;
      type_cast_2589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2589_inst_req_1;
      type_cast_2589_inst_ack_1<= rack(0);
      type_cast_2589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2701,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2589_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2599_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2599_inst_req_0;
      type_cast_2599_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2599_inst_req_1;
      type_cast_2599_inst_ack_1<= rack(0);
      type_cast_2599_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2599_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10100_2600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2619_inst
    process(sext103_2616) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2616(31 downto 0);
      type_cast_2619_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2624_inst
    process(ASHR_i32_i32_2623_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2623_wire(31 downto 0);
      shr_2625 <= tmp_var; -- 
    end process;
    type_cast_2629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2629_inst_req_0;
      type_cast_2629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2629_inst_req_1;
      type_cast_2629_inst_ack_1<= rack(0);
      type_cast_2629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2629_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2628_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2630,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2650_inst
    process(sext104_2647) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext104_2647(31 downto 0);
      type_cast_2650_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2655_inst
    process(ASHR_i32_i32_2654_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2654_wire(31 downto 0);
      shr61_2656 <= tmp_var; -- 
    end process;
    type_cast_2660_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2660_inst_req_0;
      type_cast_2660_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2660_inst_req_1;
      type_cast_2660_inst_ack_1<= rack(0);
      type_cast_2660_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2660_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2659_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom62_2661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2676_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2676_inst_req_0;
      type_cast_2676_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2676_inst_req_1;
      type_cast_2676_inst_ack_1<= rack(0);
      type_cast_2676_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2676_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2675_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_2677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2713_inst_req_0;
      type_cast_2713_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2713_inst_req_1;
      type_cast_2713_inst_ack_1<= rack(0);
      type_cast_2713_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2713_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2712_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2714,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2722_inst_req_0;
      type_cast_2722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2722_inst_req_1;
      type_cast_2722_inst_ack_1<= rack(0);
      type_cast_2722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp79_2719,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc83_2723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2739_inst_req_0;
      type_cast_2739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2739_inst_req_1;
      type_cast_2739_inst_ack_1<= rack(0);
      type_cast_2739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2738_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2740,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2391_gather_scatter
    process(LOAD_padding_2391_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2391_data_0;
      ov(15 downto 0) := iv;
      tmp27_2392 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2635_index_1_rename
    process(R_idxprom_2634_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2634_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2634_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2635_index_1_resize
    process(idxprom_2630) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2630;
      ov := iv(13 downto 0);
      R_idxprom_2634_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2635_root_address_inst
    process(array_obj_ref_2635_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2635_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2635_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2666_index_1_rename
    process(R_idxprom62_2665_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom62_2665_resized;
      ov(13 downto 0) := iv;
      R_idxprom62_2665_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2666_index_1_resize
    process(idxprom62_2661) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom62_2661;
      ov := iv(13 downto 0);
      R_idxprom62_2665_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2666_root_address_inst
    process(array_obj_ref_2666_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2666_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2666_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2328_addr_0
    process(ptr_deref_2328_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2328_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2328_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2328_base_resize
    process(iNsTr_2_2325) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2325;
      ov := iv(6 downto 0);
      ptr_deref_2328_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2328_gather_scatter
    process(ptr_deref_2328_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2328_data_0;
      ov(31 downto 0) := iv;
      tmp_2329 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2328_root_address_inst
    process(ptr_deref_2328_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2328_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2328_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2350_addr_0
    process(ptr_deref_2350_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2350_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2350_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2350_base_resize
    process(iNsTr_3_2347) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2347;
      ov := iv(6 downto 0);
      ptr_deref_2350_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2350_gather_scatter
    process(ptr_deref_2350_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2350_data_0;
      ov(31 downto 0) := iv;
      tmp11_2351 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2350_root_address_inst
    process(ptr_deref_2350_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2350_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2350_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2362_addr_0
    process(ptr_deref_2362_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2362_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2362_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2362_base_resize
    process(iNsTr_4_2359) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2359;
      ov := iv(6 downto 0);
      ptr_deref_2362_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2362_gather_scatter
    process(ptr_deref_2362_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2362_data_0;
      ov(31 downto 0) := iv;
      tmp14_2363 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2362_root_address_inst
    process(ptr_deref_2362_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2362_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2362_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2372_addr_0
    process(ptr_deref_2372_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2372_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2372_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2372_base_resize
    process(iNsTr_5_2369) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2369;
      ov := iv(0 downto 0);
      ptr_deref_2372_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2372_gather_scatter
    process(ptr_deref_2372_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2372_data_0;
      ov(15 downto 0) := iv;
      tmp22_2373 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2372_root_address_inst
    process(ptr_deref_2372_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2372_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2372_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2388_addr_0
    process(ptr_deref_2388_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2388_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2388_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2388_base_resize
    process(iNsTr_6_2385) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2385;
      ov := iv(6 downto 0);
      ptr_deref_2388_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2388_gather_scatter
    process(ptr_deref_2388_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2388_data_0;
      ov(31 downto 0) := iv;
      tmp25_2389 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2388_root_address_inst
    process(ptr_deref_2388_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2388_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2388_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2405_addr_0
    process(ptr_deref_2405_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2405_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2405_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2405_base_resize
    process(iNsTr_7_2402) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2402;
      ov := iv(0 downto 0);
      ptr_deref_2405_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2405_gather_scatter
    process(ptr_deref_2405_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2405_data_0;
      ov(15 downto 0) := iv;
      tmp33_2406 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2405_root_address_inst
    process(ptr_deref_2405_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2405_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2405_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2421_addr_0
    process(ptr_deref_2421_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2421_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2421_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2421_base_resize
    process(iNsTr_8_2418) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2418;
      ov := iv(6 downto 0);
      ptr_deref_2421_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2421_gather_scatter
    process(ptr_deref_2421_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2421_data_0;
      ov(31 downto 0) := iv;
      tmp36_2422 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2421_root_address_inst
    process(ptr_deref_2421_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2421_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2421_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2433_addr_0
    process(ptr_deref_2433_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2433_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2433_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2433_base_resize
    process(iNsTr_9_2430) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2430;
      ov := iv(6 downto 0);
      ptr_deref_2433_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2433_gather_scatter
    process(ptr_deref_2433_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2433_data_0;
      ov(31 downto 0) := iv;
      tmp45_2434 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2433_root_address_inst
    process(ptr_deref_2433_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2433_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2433_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2445_addr_0
    process(ptr_deref_2445_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2445_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2445_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2445_base_resize
    process(iNsTr_10_2442) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2442;
      ov := iv(6 downto 0);
      ptr_deref_2445_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2445_gather_scatter
    process(ptr_deref_2445_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2445_data_0;
      ov(31 downto 0) := iv;
      tmp48_2446 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2445_root_address_inst
    process(ptr_deref_2445_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2445_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2445_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2640_addr_0
    process(ptr_deref_2640_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2640_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2640_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2640_base_resize
    process(arrayidx_2637) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2637;
      ov := iv(13 downto 0);
      ptr_deref_2640_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2640_gather_scatter
    process(ptr_deref_2640_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2640_data_0;
      ov(63 downto 0) := iv;
      tmp58_2641 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2640_root_address_inst
    process(ptr_deref_2640_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2640_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2640_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2670_addr_0
    process(ptr_deref_2670_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2670_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2670_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2670_base_resize
    process(arrayidx63_2668) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx63_2668;
      ov := iv(13 downto 0);
      ptr_deref_2670_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2670_gather_scatter
    process(tmp58_2641) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp58_2641;
      ov(63 downto 0) := iv;
      ptr_deref_2670_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2670_root_address_inst
    process(ptr_deref_2670_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2670_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2670_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2689_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2688;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2689_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2689_branch_req_0,
          ack0 => if_stmt_2689_branch_ack_0,
          ack1 => if_stmt_2689_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2746_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp87_2745;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2746_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2746_branch_req_0,
          ack0 => if_stmt_2746_branch_ack_0,
          ack1 => if_stmt_2746_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2700_inst
    process(indvar_2583) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2583, type_cast_2699_wire_constant, tmp_var);
      indvarx_xnext_2701 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2708_inst
    process(input_dim1x_x1x_xph_2455) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2455, type_cast_2707_wire_constant, tmp_var);
      inc_2709 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2727_inst
    process(inc83_2723, input_dim0x_x2x_xph_2462) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc83_2723, input_dim0x_x2x_xph_2462, tmp_var);
      inc83x_xinput_dim0x_x2_2728 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2487_inst
    process(mul_2483, conv13_2473) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2483, conv13_2473, tmp_var);
      add_2488 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2502_inst
    process(mul24_2498, tmp25_2389) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul24_2498, tmp25_2389, tmp_var);
      add26_2503 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2517_inst
    process(mul35_2513, tmp36_2422) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul35_2513, tmp36_2422, tmp_var);
      add37_2518 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2534_inst
    process(sub41_2529) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub41_2529, type_cast_2533_wire_constant, tmp_var);
      sext_2535 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2555_inst
    process(sub29_2550) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub29_2550, type_cast_2554_wire_constant, tmp_var);
      sext101_2556 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2574_inst
    process(conv47_2544, mul51_2570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv47_2544, mul51_2570, tmp_var);
      add52_2575 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2604_inst
    process(mul17_2493, conv10100_2600) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul17_2493, conv10100_2600, tmp_var);
      add18_2605 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2609_inst
    process(mul53_2580, conv10100_2600) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul53_2580, conv10100_2600, tmp_var);
      add54_2610 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2682_inst
    process(conv66_2677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv66_2677, type_cast_2681_wire_constant, tmp_var);
      add67_2683 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2542_inst
    process(type_cast_2538_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2538_wire, type_cast_2541_wire_constant, tmp_var);
      ASHR_i32_i32_2542_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2563_inst
    process(type_cast_2559_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2559_wire, type_cast_2562_wire_constant, tmp_var);
      ASHR_i32_i32_2563_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2623_inst
    process(type_cast_2619_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2619_wire, type_cast_2622_wire_constant, tmp_var);
      ASHR_i32_i32_2623_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2654_inst
    process(type_cast_2650_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2650_wire, type_cast_2653_wire_constant, tmp_var);
      ASHR_i32_i32_2654_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2718_inst
    process(conv76_2714, div78_2452) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv76_2714, div78_2452, tmp_var);
      cmp79_2719 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2744_inst
    process(conv85_2740, tmp_2329) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv85_2740, tmp_2329, tmp_var);
      cmp87_2745 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2334_inst
    process(tmp_2329) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2329, type_cast_2333_wire_constant, tmp_var);
      div_2335 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2451_inst
    process(tmp14_2363) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_2363, type_cast_2450_wire_constant, tmp_var);
      div78_2452 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2595_inst
    process(indvar_2583) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2583, type_cast_2594_wire_constant, tmp_var);
      input_dim2x_x1_2596 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2482_inst
    process(tmp14_2363, conv16_2478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_2363, conv16_2478, tmp_var);
      mul_2483 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2492_inst
    process(add_2488, tmp11_2351) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2488, tmp11_2351, tmp_var);
      mul17_2493 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2497_inst
    process(conv23_2377, conv16_2478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv23_2377, conv16_2478, tmp_var);
      mul24_2498 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2512_inst
    process(conv34_2410, conv13_2473) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv34_2410, conv13_2473, tmp_var);
      mul35_2513 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2569_inst
    process(tmp48_2446, conv50_2565) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_2446, conv50_2565, tmp_var);
      mul51_2570 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2579_inst
    process(add52_2575, tmp45_2434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add52_2575, tmp45_2434, tmp_var);
      mul53_2580 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2528_inst
    process(sub40_2523) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub40_2523, type_cast_2527_wire_constant, tmp_var);
      sub41_2529 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2549_inst
    process(sub_2508) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2508, type_cast_2548_wire_constant, tmp_var);
      sub29_2550 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2615_inst
    process(add18_2605) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add18_2605, type_cast_2614_wire_constant, tmp_var);
      sext103_2616 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2646_inst
    process(add54_2610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add54_2610, type_cast_2645_wire_constant, tmp_var);
      sext104_2647 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2507_inst
    process(add26_2503, conv28_2396) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add26_2503, conv28_2396, tmp_var);
      sub_2508 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2522_inst
    process(add37_2518, conv28_2396) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add37_2518, conv28_2396, tmp_var);
      sub40_2523 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2687_inst
    process(add67_2683, tmp11_2351) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add67_2683, tmp11_2351, tmp_var);
      cmp_2688 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_2635_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2634_scaled;
      array_obj_ref_2635_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2635_index_offset_req_0;
      array_obj_ref_2635_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2635_index_offset_req_1;
      array_obj_ref_2635_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_2666_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom62_2665_scaled;
      array_obj_ref_2666_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2666_index_offset_req_0;
      array_obj_ref_2666_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2666_index_offset_req_1;
      array_obj_ref_2666_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_2471_inst
    process(input_dim1x_x1x_xph_2455) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2455, tmp_var);
      type_cast_2471_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2476_inst
    process(input_dim0x_x2x_xph_2462) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2462, tmp_var);
      type_cast_2476_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2628_inst
    process(shr_2625) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2625, tmp_var);
      type_cast_2628_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2659_inst
    process(shr61_2656) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr61_2656, tmp_var);
      type_cast_2659_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2675_inst
    process(input_dim2x_x1_2596) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2596, tmp_var);
      type_cast_2675_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2712_inst
    process(inc_2709) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2709, tmp_var);
      type_cast_2712_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2738_inst
    process(inc83x_xinput_dim0x_x2_2728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc83x_xinput_dim0x_x2_2728, tmp_var);
      type_cast_2738_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2391_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2391_load_0_req_0;
      LOAD_padding_2391_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2391_load_0_req_1;
      LOAD_padding_2391_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2391_word_address_0;
      LOAD_padding_2391_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2362_load_0 ptr_deref_2350_load_0 ptr_deref_2328_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2362_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2350_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2328_load_0_req_0;
      ptr_deref_2362_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2350_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2328_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2362_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2350_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2328_load_0_req_1;
      ptr_deref_2362_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2350_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2328_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2362_word_address_0 & ptr_deref_2350_word_address_0 & ptr_deref_2328_word_address_0;
      ptr_deref_2362_data_0 <= data_out(95 downto 64);
      ptr_deref_2350_data_0 <= data_out(63 downto 32);
      ptr_deref_2328_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2372_load_0 ptr_deref_2405_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2372_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2405_load_0_req_0;
      ptr_deref_2372_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2405_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2372_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2405_load_0_req_1;
      ptr_deref_2372_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2405_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2372_word_address_0 & ptr_deref_2405_word_address_0;
      ptr_deref_2372_data_0 <= data_out(31 downto 16);
      ptr_deref_2405_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2421_load_0 ptr_deref_2388_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2421_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2388_load_0_req_0;
      ptr_deref_2421_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2388_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2421_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2388_load_0_req_1;
      ptr_deref_2421_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2388_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2421_word_address_0 & ptr_deref_2388_word_address_0;
      ptr_deref_2421_data_0 <= data_out(63 downto 32);
      ptr_deref_2388_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2445_load_0 ptr_deref_2433_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2445_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2433_load_0_req_0;
      ptr_deref_2445_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2433_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2445_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2433_load_0_req_1;
      ptr_deref_2445_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2433_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2445_word_address_0 & ptr_deref_2433_word_address_0;
      ptr_deref_2445_data_0 <= data_out(63 downto 32);
      ptr_deref_2433_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2640_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2640_load_0_req_0;
      ptr_deref_2640_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2640_load_0_req_1;
      ptr_deref_2640_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2640_word_address_0;
      ptr_deref_2640_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2670_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2670_store_0_req_0;
      ptr_deref_2670_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2670_store_0_req_1;
      ptr_deref_2670_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2670_word_address_0;
      data_in <= ptr_deref_2670_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2315_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_start_2315_inst_req_0;
      RPIPE_Block2_start_2315_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_start_2315_inst_req_1;
      RPIPE_Block2_start_2315_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2316 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2754_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2754_inst_req_0;
      WPIPE_Block2_done_2754_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2754_inst_req_1;
      WPIPE_Block2_done_2754_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2316;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_7773_start: Boolean;
  signal convTransposeD_CP_7773_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2809_inst_req_0 : boolean;
  signal type_cast_2809_inst_ack_0 : boolean;
  signal ptr_deref_2799_load_0_req_0 : boolean;
  signal type_cast_2787_inst_ack_1 : boolean;
  signal LOAD_padding_2850_load_0_ack_1 : boolean;
  signal LOAD_padding_2850_load_0_req_0 : boolean;
  signal LOAD_padding_2850_load_0_ack_0 : boolean;
  signal LOAD_padding_2850_load_0_req_1 : boolean;
  signal ptr_deref_2847_load_0_ack_1 : boolean;
  signal type_cast_2809_inst_req_1 : boolean;
  signal type_cast_2854_inst_ack_0 : boolean;
  signal type_cast_2854_inst_req_1 : boolean;
  signal type_cast_2854_inst_req_0 : boolean;
  signal type_cast_2809_inst_ack_1 : boolean;
  signal ptr_deref_2799_load_0_ack_1 : boolean;
  signal ptr_deref_2831_load_0_ack_1 : boolean;
  signal ptr_deref_2847_load_0_req_0 : boolean;
  signal ptr_deref_2847_load_0_ack_0 : boolean;
  signal ptr_deref_2821_load_0_req_1 : boolean;
  signal ptr_deref_2821_load_0_ack_1 : boolean;
  signal ptr_deref_2847_load_0_req_1 : boolean;
  signal ptr_deref_2831_load_0_req_1 : boolean;
  signal type_cast_2835_inst_req_0 : boolean;
  signal type_cast_2835_inst_ack_0 : boolean;
  signal type_cast_2835_inst_req_1 : boolean;
  signal type_cast_2787_inst_req_1 : boolean;
  signal type_cast_2835_inst_ack_1 : boolean;
  signal ptr_deref_2831_load_0_req_0 : boolean;
  signal ptr_deref_2831_load_0_ack_0 : boolean;
  signal ptr_deref_2821_load_0_req_0 : boolean;
  signal ptr_deref_2821_load_0_ack_0 : boolean;
  signal type_cast_2868_inst_req_0 : boolean;
  signal type_cast_2868_inst_ack_0 : boolean;
  signal ptr_deref_2864_load_0_req_0 : boolean;
  signal type_cast_2854_inst_ack_1 : boolean;
  signal ptr_deref_2864_load_0_ack_0 : boolean;
  signal ptr_deref_2799_load_0_req_1 : boolean;
  signal type_cast_2868_inst_req_1 : boolean;
  signal type_cast_2868_inst_ack_1 : boolean;
  signal ptr_deref_2799_load_0_ack_0 : boolean;
  signal ptr_deref_2864_load_0_req_1 : boolean;
  signal ptr_deref_2864_load_0_ack_1 : boolean;
  signal ptr_deref_2880_load_0_req_0 : boolean;
  signal ptr_deref_2880_load_0_ack_0 : boolean;
  signal ptr_deref_2880_load_0_req_1 : boolean;
  signal ptr_deref_2880_load_0_ack_1 : boolean;
  signal type_cast_2787_inst_ack_0 : boolean;
  signal type_cast_2787_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2764_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2764_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2764_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2764_inst_ack_1 : boolean;
  signal ptr_deref_2777_load_0_req_0 : boolean;
  signal ptr_deref_2777_load_0_ack_0 : boolean;
  signal ptr_deref_2777_load_0_req_1 : boolean;
  signal ptr_deref_2777_load_0_ack_1 : boolean;
  signal ptr_deref_2892_load_0_req_0 : boolean;
  signal ptr_deref_2892_load_0_ack_0 : boolean;
  signal ptr_deref_2892_load_0_req_1 : boolean;
  signal ptr_deref_2892_load_0_ack_1 : boolean;
  signal ptr_deref_2904_load_0_req_0 : boolean;
  signal ptr_deref_2904_load_0_ack_0 : boolean;
  signal ptr_deref_2904_load_0_req_1 : boolean;
  signal ptr_deref_2904_load_0_ack_1 : boolean;
  signal type_cast_2924_inst_req_0 : boolean;
  signal type_cast_2924_inst_ack_0 : boolean;
  signal type_cast_2924_inst_req_1 : boolean;
  signal type_cast_2924_inst_ack_1 : boolean;
  signal type_cast_2929_inst_req_0 : boolean;
  signal type_cast_2929_inst_ack_0 : boolean;
  signal type_cast_2929_inst_req_1 : boolean;
  signal type_cast_2929_inst_ack_1 : boolean;
  signal type_cast_3051_inst_req_0 : boolean;
  signal type_cast_3051_inst_ack_0 : boolean;
  signal type_cast_3051_inst_req_1 : boolean;
  signal type_cast_3051_inst_ack_1 : boolean;
  signal type_cast_3081_inst_req_0 : boolean;
  signal type_cast_3081_inst_ack_0 : boolean;
  signal type_cast_3081_inst_req_1 : boolean;
  signal type_cast_3081_inst_ack_1 : boolean;
  signal array_obj_ref_3087_index_offset_req_0 : boolean;
  signal array_obj_ref_3087_index_offset_ack_0 : boolean;
  signal array_obj_ref_3087_index_offset_req_1 : boolean;
  signal array_obj_ref_3087_index_offset_ack_1 : boolean;
  signal addr_of_3088_final_reg_req_0 : boolean;
  signal addr_of_3088_final_reg_ack_0 : boolean;
  signal addr_of_3088_final_reg_req_1 : boolean;
  signal addr_of_3088_final_reg_ack_1 : boolean;
  signal ptr_deref_3092_load_0_req_0 : boolean;
  signal ptr_deref_3092_load_0_ack_0 : boolean;
  signal ptr_deref_3092_load_0_req_1 : boolean;
  signal ptr_deref_3092_load_0_ack_1 : boolean;
  signal type_cast_3112_inst_req_0 : boolean;
  signal type_cast_3112_inst_ack_0 : boolean;
  signal type_cast_3112_inst_req_1 : boolean;
  signal type_cast_3112_inst_ack_1 : boolean;
  signal array_obj_ref_3118_index_offset_req_0 : boolean;
  signal array_obj_ref_3118_index_offset_ack_0 : boolean;
  signal array_obj_ref_3118_index_offset_req_1 : boolean;
  signal array_obj_ref_3118_index_offset_ack_1 : boolean;
  signal addr_of_3119_final_reg_req_0 : boolean;
  signal addr_of_3119_final_reg_ack_0 : boolean;
  signal addr_of_3119_final_reg_req_1 : boolean;
  signal addr_of_3119_final_reg_ack_1 : boolean;
  signal ptr_deref_3122_store_0_req_0 : boolean;
  signal ptr_deref_3122_store_0_ack_0 : boolean;
  signal ptr_deref_3122_store_0_req_1 : boolean;
  signal ptr_deref_3122_store_0_ack_1 : boolean;
  signal type_cast_3128_inst_req_0 : boolean;
  signal type_cast_3128_inst_ack_0 : boolean;
  signal type_cast_3128_inst_req_1 : boolean;
  signal type_cast_3128_inst_ack_1 : boolean;
  signal if_stmt_3141_branch_req_0 : boolean;
  signal if_stmt_3141_branch_ack_1 : boolean;
  signal if_stmt_3141_branch_ack_0 : boolean;
  signal type_cast_3165_inst_req_0 : boolean;
  signal type_cast_3165_inst_ack_0 : boolean;
  signal type_cast_3165_inst_req_1 : boolean;
  signal type_cast_3165_inst_ack_1 : boolean;
  signal if_stmt_3172_branch_req_0 : boolean;
  signal if_stmt_3172_branch_ack_1 : boolean;
  signal if_stmt_3172_branch_ack_0 : boolean;
  signal type_cast_3193_inst_req_0 : boolean;
  signal type_cast_3193_inst_ack_0 : boolean;
  signal type_cast_3193_inst_req_1 : boolean;
  signal type_cast_3193_inst_ack_1 : boolean;
  signal type_cast_3213_inst_req_0 : boolean;
  signal type_cast_3213_inst_ack_0 : boolean;
  signal type_cast_3213_inst_req_1 : boolean;
  signal type_cast_3213_inst_ack_1 : boolean;
  signal if_stmt_3220_branch_req_0 : boolean;
  signal if_stmt_3220_branch_ack_1 : boolean;
  signal if_stmt_3220_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_3228_inst_req_0 : boolean;
  signal WPIPE_Block3_done_3228_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_3228_inst_req_1 : boolean;
  signal WPIPE_Block3_done_3228_inst_ack_1 : boolean;
  signal type_cast_2911_inst_req_0 : boolean;
  signal type_cast_2911_inst_ack_0 : boolean;
  signal type_cast_2911_inst_req_1 : boolean;
  signal type_cast_2911_inst_ack_1 : boolean;
  signal phi_stmt_2908_req_0 : boolean;
  signal type_cast_2917_inst_req_0 : boolean;
  signal type_cast_2917_inst_ack_0 : boolean;
  signal type_cast_2917_inst_req_1 : boolean;
  signal type_cast_2917_inst_ack_1 : boolean;
  signal phi_stmt_2914_req_0 : boolean;
  signal type_cast_2913_inst_req_0 : boolean;
  signal type_cast_2913_inst_ack_0 : boolean;
  signal type_cast_2913_inst_req_1 : boolean;
  signal type_cast_2913_inst_ack_1 : boolean;
  signal phi_stmt_2908_req_1 : boolean;
  signal type_cast_2919_inst_req_0 : boolean;
  signal type_cast_2919_inst_ack_0 : boolean;
  signal type_cast_2919_inst_req_1 : boolean;
  signal type_cast_2919_inst_ack_1 : boolean;
  signal phi_stmt_2914_req_1 : boolean;
  signal phi_stmt_2908_ack_0 : boolean;
  signal phi_stmt_2914_ack_0 : boolean;
  signal type_cast_3041_inst_req_0 : boolean;
  signal type_cast_3041_inst_ack_0 : boolean;
  signal type_cast_3041_inst_req_1 : boolean;
  signal type_cast_3041_inst_ack_1 : boolean;
  signal phi_stmt_3035_req_1 : boolean;
  signal phi_stmt_3035_req_0 : boolean;
  signal phi_stmt_3035_ack_0 : boolean;
  signal type_cast_3206_inst_req_0 : boolean;
  signal type_cast_3206_inst_ack_0 : boolean;
  signal type_cast_3206_inst_req_1 : boolean;
  signal type_cast_3206_inst_ack_1 : boolean;
  signal phi_stmt_3203_req_0 : boolean;
  signal type_cast_3200_inst_req_0 : boolean;
  signal type_cast_3200_inst_ack_0 : boolean;
  signal type_cast_3200_inst_req_1 : boolean;
  signal type_cast_3200_inst_ack_1 : boolean;
  signal phi_stmt_3197_req_0 : boolean;
  signal type_cast_3208_inst_req_0 : boolean;
  signal type_cast_3208_inst_ack_0 : boolean;
  signal type_cast_3208_inst_req_1 : boolean;
  signal type_cast_3208_inst_ack_1 : boolean;
  signal phi_stmt_3203_req_1 : boolean;
  signal type_cast_3202_inst_req_0 : boolean;
  signal type_cast_3202_inst_ack_0 : boolean;
  signal type_cast_3202_inst_req_1 : boolean;
  signal type_cast_3202_inst_ack_1 : boolean;
  signal phi_stmt_3197_req_1 : boolean;
  signal phi_stmt_3197_ack_0 : boolean;
  signal phi_stmt_3203_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_7773_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7773_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_7773_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7773_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_7773: Block -- control-path 
    signal convTransposeD_CP_7773_elements: BooleanArray(116 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_7773_elements(0) <= convTransposeD_CP_7773_start;
    convTransposeD_CP_7773_symbol <= convTransposeD_CP_7773_elements(74);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2762/$entry
      -- CP-element group 0: 	 branch_block_stmt_2762/branch_block_stmt_2762__entry__
      -- CP-element group 0: 	 branch_block_stmt_2762/assign_stmt_2765__entry__
      -- CP-element group 0: 	 branch_block_stmt_2762/assign_stmt_2765/$entry
      -- CP-element group 0: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_Sample/rr
      -- 
    rr_7831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(0), ack => RPIPE_Block3_start_2764_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_Update/cr
      -- 
    ra_7832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2764_inst_ack_0, ack => convTransposeD_CP_7773_elements(1)); -- 
    cr_7836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(1), ack => RPIPE_Block3_start_2764_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	31 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	32 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (268) 
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2765__exit__
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905__entry__
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2765/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2765/RPIPE_Block3_start_2764_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/word_access_complete/word_0/cr
      -- 
    ca_7837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2764_inst_ack_1, ack => convTransposeD_CP_7773_elements(2)); -- 
    rr_7937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2799_load_0_req_0); -- 
    rr_8148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => LOAD_padding_2850_load_0_req_0); -- 
    cr_8159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => LOAD_padding_2850_load_0_req_1); -- 
    cr_7967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => type_cast_2809_inst_req_1); -- 
    cr_8178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => type_cast_2854_inst_req_1); -- 
    rr_8115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2847_load_0_req_0); -- 
    cr_8012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2821_load_0_req_1); -- 
    cr_8126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2847_load_0_req_1); -- 
    cr_8062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2831_load_0_req_1); -- 
    cr_8081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => type_cast_2835_inst_req_1); -- 
    cr_7903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => type_cast_2787_inst_req_1); -- 
    rr_8051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2831_load_0_req_0); -- 
    rr_8001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2821_load_0_req_0); -- 
    rr_8212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2864_load_0_req_0); -- 
    cr_7948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2799_load_0_req_1); -- 
    cr_8242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => type_cast_2868_inst_req_1); -- 
    cr_8223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2864_load_0_req_1); -- 
    rr_8276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2880_load_0_req_0); -- 
    cr_8287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2880_load_0_req_1); -- 
    rr_7873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2777_load_0_req_0); -- 
    cr_7884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2777_load_0_req_1); -- 
    rr_8326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2892_load_0_req_0); -- 
    cr_8337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2892_load_0_req_1); -- 
    rr_8376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2904_load_0_req_0); -- 
    cr_8387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(2), ack => ptr_deref_2904_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Sample/word_access_start/word_0/ra
      -- 
    ra_7874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2777_load_0_ack_0, ack => convTransposeD_CP_7773_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/ptr_deref_2777_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/ptr_deref_2777_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/ptr_deref_2777_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/ptr_deref_2777_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2777_Update/word_access_complete/word_0/ca
      -- 
    ca_7885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2777_load_0_ack_1, ack => convTransposeD_CP_7773_elements(4)); -- 
    rr_7898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(4), ack => type_cast_2787_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_Sample/ra
      -- 
    ra_7899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2787_inst_ack_0, ack => convTransposeD_CP_7773_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	33 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2787_Update/$exit
      -- 
    ca_7904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2787_inst_ack_1, ack => convTransposeD_CP_7773_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Sample/word_access_start/word_0/ra
      -- 
    ra_7938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2799_load_0_ack_0, ack => convTransposeD_CP_7773_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/ptr_deref_2799_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/ptr_deref_2799_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/ptr_deref_2799_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2799_Update/ptr_deref_2799_Merge/$exit
      -- 
    ca_7949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2799_load_0_ack_1, ack => convTransposeD_CP_7773_elements(8)); -- 
    rr_7962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(8), ack => type_cast_2809_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_sample_completed_
      -- 
    ra_7963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2809_inst_ack_0, ack => convTransposeD_CP_7773_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	33 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2809_Update/ca
      -- 
    ca_7968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2809_inst_ack_1, ack => convTransposeD_CP_7773_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Sample/word_access_start/word_0/ra
      -- 
    ra_8002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2821_load_0_ack_0, ack => convTransposeD_CP_7773_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	33 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/ptr_deref_2821_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/ptr_deref_2821_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/ptr_deref_2821_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_Update/ptr_deref_2821_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2821_update_completed_
      -- 
    ca_8013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2821_load_0_ack_1, ack => convTransposeD_CP_7773_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Sample/$exit
      -- 
    ra_8052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2831_load_0_ack_0, ack => convTransposeD_CP_7773_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/ptr_deref_2831_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/ptr_deref_2831_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/ptr_deref_2831_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/ptr_deref_2831_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2831_update_completed_
      -- 
    ca_8063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2831_load_0_ack_1, ack => convTransposeD_CP_7773_elements(14)); -- 
    rr_8076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(14), ack => type_cast_2835_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_sample_completed_
      -- 
    ra_8077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2835_inst_ack_0, ack => convTransposeD_CP_7773_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	33 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2835_Update/ca
      -- 
    ca_8082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2835_inst_ack_1, ack => convTransposeD_CP_7773_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Sample/word_access_start/word_0/ra
      -- CP-element group 17: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Sample/$exit
      -- 
    ra_8116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2847_load_0_ack_0, ack => convTransposeD_CP_7773_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/ptr_deref_2847_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/ptr_deref_2847_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/ptr_deref_2847_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2847_Update/ptr_deref_2847_Merge/merge_ack
      -- 
    ca_8127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2847_load_0_ack_1, ack => convTransposeD_CP_7773_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Sample/word_access_start/word_0/ra
      -- 
    ra_8149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2850_load_0_ack_0, ack => convTransposeD_CP_7773_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/LOAD_padding_2850_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/LOAD_padding_2850_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/LOAD_padding_2850_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/LOAD_padding_2850_Update/LOAD_padding_2850_Merge/$entry
      -- 
    ca_8160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2850_load_0_ack_1, ack => convTransposeD_CP_7773_elements(20)); -- 
    rr_8173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(20), ack => type_cast_2854_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_sample_completed_
      -- 
    ra_8174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2854_inst_ack_0, ack => convTransposeD_CP_7773_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	33 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2854_Update/ca
      -- 
    ca_8179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2854_inst_ack_1, ack => convTransposeD_CP_7773_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Sample/word_access_start/word_0/ra
      -- 
    ra_8213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2864_load_0_ack_0, ack => convTransposeD_CP_7773_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (12) 
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/ptr_deref_2864_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/ptr_deref_2864_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/ptr_deref_2864_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2864_Update/ptr_deref_2864_Merge/$entry
      -- 
    ca_8224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2864_load_0_ack_1, ack => convTransposeD_CP_7773_elements(24)); -- 
    rr_8237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(24), ack => type_cast_2868_inst_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_sample_completed_
      -- 
    ra_8238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2868_inst_ack_0, ack => convTransposeD_CP_7773_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	33 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/type_cast_2868_Update/ca
      -- 
    ca_8243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2868_inst_ack_1, ack => convTransposeD_CP_7773_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Sample/word_access_start/word_0/ra
      -- 
    ra_8277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2880_load_0_ack_0, ack => convTransposeD_CP_7773_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	33 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/ptr_deref_2880_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/ptr_deref_2880_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/ptr_deref_2880_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2880_Update/ptr_deref_2880_Merge/merge_ack
      -- 
    ca_8288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2880_load_0_ack_1, ack => convTransposeD_CP_7773_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Sample/word_access_start/word_0/ra
      -- 
    ra_8327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_load_0_ack_0, ack => convTransposeD_CP_7773_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/ptr_deref_2892_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/ptr_deref_2892_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/ptr_deref_2892_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2892_Update/ptr_deref_2892_Merge/merge_ack
      -- 
    ca_8338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_load_0_ack_1, ack => convTransposeD_CP_7773_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	2 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Sample/word_access_start/word_0/ra
      -- 
    ra_8377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_0_ack_0, ack => convTransposeD_CP_7773_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/ptr_deref_2904_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/ptr_deref_2904_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/ptr_deref_2904_Merge/merge_req
      -- CP-element group 32: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/ptr_deref_2904_Update/ptr_deref_2904_Merge/merge_ack
      -- 
    ca_8388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_0_ack_1, ack => convTransposeD_CP_7773_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  place  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	12 
    -- CP-element group 33: 	6 
    -- CP-element group 33: 	18 
    -- CP-element group 33: 	10 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	30 
    -- CP-element group 33: 	26 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	75 
    -- CP-element group 33: 	76 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	79 
    -- CP-element group 33:  members (20) 
      -- CP-element group 33: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905__exit__
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter
      -- CP-element group 33: 	 branch_block_stmt_2762/assign_stmt_2774_to_assign_stmt_2905/$exit
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Update/cr
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/cr
      -- 
    rr_8822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(33), ack => type_cast_2911_inst_req_0); -- 
    cr_8827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(33), ack => type_cast_2911_inst_req_1); -- 
    rr_8845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(33), ack => type_cast_2917_inst_req_0); -- 
    cr_8850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(33), ack => type_cast_2917_inst_req_1); -- 
    convTransposeD_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(12) & convTransposeD_CP_7773_elements(6) & convTransposeD_CP_7773_elements(18) & convTransposeD_CP_7773_elements(10) & convTransposeD_CP_7773_elements(22) & convTransposeD_CP_7773_elements(28) & convTransposeD_CP_7773_elements(16) & convTransposeD_CP_7773_elements(30) & convTransposeD_CP_7773_elements(26) & convTransposeD_CP_7773_elements(32);
      gj_convTransposeD_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	92 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_Sample/ra
      -- 
    ra_8405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2924_inst_ack_0, ack => convTransposeD_CP_7773_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	92 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_Update/ca
      -- 
    ca_8410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2924_inst_ack_1, ack => convTransposeD_CP_7773_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	92 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_Sample/ra
      -- 
    ra_8419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2929_inst_ack_0, ack => convTransposeD_CP_7773_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_Update/ca
      -- 
    ca_8424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2929_inst_ack_1, ack => convTransposeD_CP_7773_elements(37)); -- 
    -- CP-element group 38:  join  transition  place  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	96 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032__exit__
      -- CP-element group 38: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 38: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/$exit
      -- CP-element group 38: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3035/$entry
      -- CP-element group 38: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/$entry
      -- 
    convTransposeD_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(37) & convTransposeD_CP_7773_elements(35);
      gj_convTransposeD_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	98 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_Sample/ra
      -- 
    ra_8436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3051_inst_ack_0, ack => convTransposeD_CP_7773_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	98 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_Sample/rr
      -- 
    ca_8441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3051_inst_ack_1, ack => convTransposeD_CP_7773_elements(40)); -- 
    rr_8559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(40), ack => type_cast_3112_inst_req_0); -- 
    rr_8449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(40), ack => type_cast_3081_inst_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_Sample/ra
      -- 
    ra_8450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3081_inst_ack_0, ack => convTransposeD_CP_7773_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	98 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (16) 
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_resized_1
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_scaled_1
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_computed_1
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_resize_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_resize_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_resize_1/index_resize_req
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_resize_1/index_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_scale_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_scale_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_scale_1/scale_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_index_scale_1/scale_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_Sample/req
      -- 
    ca_8455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3081_inst_ack_1, ack => convTransposeD_CP_7773_elements(42)); -- 
    req_8480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(42), ack => array_obj_ref_3087_index_offset_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	60 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_sample_complete
      -- CP-element group 43: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_Sample/ack
      -- 
    ack_8481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3087_index_offset_ack_0, ack => convTransposeD_CP_7773_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	98 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (11) 
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_offset_calculated
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_Update/ack
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_request/$entry
      -- CP-element group 44: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_request/req
      -- 
    ack_8486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3087_index_offset_ack_1, ack => convTransposeD_CP_7773_elements(44)); -- 
    req_8495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(44), ack => addr_of_3088_final_reg_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_request/$exit
      -- CP-element group 45: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_request/ack
      -- 
    ack_8496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3088_final_reg_ack_0, ack => convTransposeD_CP_7773_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	98 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (24) 
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_complete/ack
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_word_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_root_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_address_resized
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_addr_resize/$entry
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_addr_resize/$exit
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_addr_resize/base_resize_req
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_addr_resize/base_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_plus_offset/$entry
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_plus_offset/$exit
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_plus_offset/sum_rename_req
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_base_plus_offset/sum_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_word_addrgen/$entry
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_word_addrgen/$exit
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_word_addrgen/root_register_req
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_word_addrgen/root_register_ack
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Sample/word_access_start/$entry
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Sample/word_access_start/word_0/$entry
      -- CP-element group 46: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Sample/word_access_start/word_0/rr
      -- 
    ack_8501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3088_final_reg_ack_1, ack => convTransposeD_CP_7773_elements(46)); -- 
    rr_8534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(46), ack => ptr_deref_3092_load_0_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Sample/word_access_start/$exit
      -- CP-element group 47: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Sample/word_access_start/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Sample/word_access_start/word_0/ra
      -- 
    ra_8535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3092_load_0_ack_0, ack => convTransposeD_CP_7773_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	98 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	55 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/word_access_complete/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/word_access_complete/word_0/ca
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/ptr_deref_3092_Merge/$entry
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/ptr_deref_3092_Merge/$exit
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/ptr_deref_3092_Merge/merge_req
      -- CP-element group 48: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/ptr_deref_3092_Merge/merge_ack
      -- 
    ca_8546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3092_load_0_ack_1, ack => convTransposeD_CP_7773_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	40 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_Sample/ra
      -- 
    ra_8560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3112_inst_ack_0, ack => convTransposeD_CP_7773_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	98 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (16) 
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_resized_1
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_scaled_1
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_computed_1
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_resize_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_resize_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_resize_1/index_resize_req
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_resize_1/index_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_scale_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_scale_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_scale_1/scale_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_index_scale_1/scale_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_Sample/req
      -- 
    ca_8565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3112_inst_ack_1, ack => convTransposeD_CP_7773_elements(50)); -- 
    req_8590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(50), ack => array_obj_ref_3118_index_offset_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	60 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_sample_complete
      -- CP-element group 51: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_Sample/ack
      -- 
    ack_8591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3118_index_offset_ack_0, ack => convTransposeD_CP_7773_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	98 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (11) 
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_offset_calculated
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_request/$entry
      -- CP-element group 52: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_request/req
      -- 
    ack_8596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3118_index_offset_ack_1, ack => convTransposeD_CP_7773_elements(52)); -- 
    req_8605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(52), ack => addr_of_3119_final_reg_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_request/$exit
      -- CP-element group 53: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_request/ack
      -- 
    ack_8606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3119_final_reg_ack_0, ack => convTransposeD_CP_7773_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	98 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (19) 
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_complete/$exit
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_complete/ack
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_word_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_root_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_address_resized
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_addr_resize/$entry
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_addr_resize/$exit
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_addr_resize/base_resize_req
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_addr_resize/base_resize_ack
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_plus_offset/$entry
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_plus_offset/$exit
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_plus_offset/sum_rename_req
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_base_plus_offset/sum_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_word_addrgen/$entry
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_word_addrgen/$exit
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_word_addrgen/root_register_req
      -- CP-element group 54: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_word_addrgen/root_register_ack
      -- 
    ack_8611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3119_final_reg_ack_1, ack => convTransposeD_CP_7773_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	48 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/ptr_deref_3122_Split/$entry
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/ptr_deref_3122_Split/$exit
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/ptr_deref_3122_Split/split_req
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/ptr_deref_3122_Split/split_ack
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/word_access_start/word_0/rr
      -- 
    rr_8649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(55), ack => ptr_deref_3122_store_0_req_0); -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(48) & convTransposeD_CP_7773_elements(54);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Sample/word_access_start/word_0/ra
      -- 
    ra_8650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3122_store_0_ack_0, ack => convTransposeD_CP_7773_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	98 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	60 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Update/word_access_complete/word_0/ca
      -- 
    ca_8661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3122_store_0_ack_1, ack => convTransposeD_CP_7773_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	98 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_Sample/ra
      -- 
    ra_8670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3128_inst_ack_0, ack => convTransposeD_CP_7773_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	98 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_Update/ca
      -- 
    ca_8675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3128_inst_ack_1, ack => convTransposeD_CP_7773_elements(59)); -- 
    -- CP-element group 60:  branch  join  transition  place  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	43 
    -- CP-element group 60: 	57 
    -- CP-element group 60: 	51 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (10) 
      -- CP-element group 60: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140__exit__
      -- CP-element group 60: 	 branch_block_stmt_2762/if_stmt_3141__entry__
      -- CP-element group 60: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/$exit
      -- CP-element group 60: 	 branch_block_stmt_2762/if_stmt_3141_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2762/if_stmt_3141_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_2762/if_stmt_3141_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_2762/if_stmt_3141_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_2762/R_cmp_3142_place
      -- CP-element group 60: 	 branch_block_stmt_2762/if_stmt_3141_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2762/if_stmt_3141_else_link/$entry
      -- 
    branch_req_8683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(60), ack => if_stmt_3141_branch_req_0); -- 
    convTransposeD_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(43) & convTransposeD_CP_7773_elements(57) & convTransposeD_CP_7773_elements(51) & convTransposeD_CP_7773_elements(59);
      gj_convTransposeD_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	93 
    -- CP-element group 61: 	94 
    -- CP-element group 61:  members (24) 
      -- CP-element group 61: 	 branch_block_stmt_2762/merge_stmt_3147__exit__
      -- CP-element group 61: 	 branch_block_stmt_2762/assign_stmt_3153__entry__
      -- CP-element group 61: 	 branch_block_stmt_2762/assign_stmt_3153__exit__
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody
      -- CP-element group 61: 	 branch_block_stmt_2762/if_stmt_3141_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_2762/if_stmt_3141_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_2762/whilex_xbody_ifx_xthen
      -- CP-element group 61: 	 branch_block_stmt_2762/assign_stmt_3153/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/assign_stmt_3153/$exit
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/Update/cr
      -- CP-element group 61: 	 branch_block_stmt_2762/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_2762/merge_stmt_3147_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_2762/merge_stmt_3147_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_2762/merge_stmt_3147_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_2762/merge_stmt_3147_PhiAck/dummy
      -- 
    if_choice_transition_8688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3141_branch_ack_1, ack => convTransposeD_CP_7773_elements(61)); -- 
    rr_8926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(61), ack => type_cast_3041_inst_req_0); -- 
    cr_8931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(61), ack => type_cast_3041_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (18) 
      -- CP-element group 62: 	 branch_block_stmt_2762/merge_stmt_3155__exit__
      -- CP-element group 62: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171__entry__
      -- CP-element group 62: 	 branch_block_stmt_2762/if_stmt_3141_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_2762/if_stmt_3141_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_2762/whilex_xbody_ifx_xelse
      -- CP-element group 62: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/$entry
      -- CP-element group 62: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_2762/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_2762/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_2762/merge_stmt_3155_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_2762/merge_stmt_3155_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_2762/merge_stmt_3155_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_2762/merge_stmt_3155_PhiAck/dummy
      -- 
    else_choice_transition_8692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3141_branch_ack_0, ack => convTransposeD_CP_7773_elements(62)); -- 
    rr_8708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(62), ack => type_cast_3165_inst_req_0); -- 
    cr_8713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(62), ack => type_cast_3165_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_Sample/ra
      -- 
    ra_8709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3165_inst_ack_0, ack => convTransposeD_CP_7773_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171__exit__
      -- CP-element group 64: 	 branch_block_stmt_2762/if_stmt_3172__entry__
      -- CP-element group 64: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/$exit
      -- CP-element group 64: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2762/assign_stmt_3161_to_assign_stmt_3171/type_cast_3165_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2762/if_stmt_3172_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2762/if_stmt_3172_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_2762/if_stmt_3172_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_2762/if_stmt_3172_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_2762/R_cmp81_3173_place
      -- CP-element group 64: 	 branch_block_stmt_2762/if_stmt_3172_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2762/if_stmt_3172_else_link/$entry
      -- 
    ca_8714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3165_inst_ack_1, ack => convTransposeD_CP_7773_elements(64)); -- 
    branch_req_8722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(64), ack => if_stmt_3172_branch_req_0); -- 
    -- CP-element group 65:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (18) 
      -- CP-element group 65: 	 branch_block_stmt_2762/merge_stmt_3178__exit__
      -- CP-element group 65: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194__entry__
      -- CP-element group 65: 	 branch_block_stmt_2762/if_stmt_3172_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2762/if_stmt_3172_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2762/ifx_xelse_ifx_xthen83
      -- CP-element group 65: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/$entry
      -- CP-element group 65: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2762/ifx_xelse_ifx_xthen83_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2762/ifx_xelse_ifx_xthen83_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_2762/merge_stmt_3178_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_2762/merge_stmt_3178_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_2762/merge_stmt_3178_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_2762/merge_stmt_3178_PhiAck/dummy
      -- 
    if_choice_transition_8727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3172_branch_ack_1, ack => convTransposeD_CP_7773_elements(65)); -- 
    rr_8744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(65), ack => type_cast_3193_inst_req_0); -- 
    cr_8749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(65), ack => type_cast_3193_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	99 
    -- CP-element group 66: 	100 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	103 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_2762/if_stmt_3172_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_2762/if_stmt_3172_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3172_branch_ack_0, ack => convTransposeD_CP_7773_elements(66)); -- 
    rr_9000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(66), ack => type_cast_3206_inst_req_0); -- 
    cr_9005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(66), ack => type_cast_3206_inst_req_1); -- 
    rr_9023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(66), ack => type_cast_3200_inst_req_0); -- 
    cr_9028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(66), ack => type_cast_3200_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_Sample/ra
      -- 
    ra_8745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3193_inst_ack_0, ack => convTransposeD_CP_7773_elements(67)); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	106 
    -- CP-element group 68: 	107 
    -- CP-element group 68: 	109 
    -- CP-element group 68: 	110 
    -- CP-element group 68:  members (23) 
      -- CP-element group 68: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194__exit__
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend
      -- CP-element group 68: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/$exit
      -- CP-element group 68: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2762/assign_stmt_3184_to_assign_stmt_3194/type_cast_3193_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/Update/cr
      -- 
    ca_8750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3193_inst_ack_1, ack => convTransposeD_CP_7773_elements(68)); -- 
    rr_9049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(68), ack => type_cast_3208_inst_req_0); -- 
    cr_9054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(68), ack => type_cast_3208_inst_req_1); -- 
    rr_9072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(68), ack => type_cast_3202_inst_req_0); -- 
    cr_9077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(68), ack => type_cast_3202_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	116 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_Sample/ra
      -- 
    ra_8762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3213_inst_ack_0, ack => convTransposeD_CP_7773_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	116 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219__exit__
      -- CP-element group 70: 	 branch_block_stmt_2762/if_stmt_3220__entry__
      -- CP-element group 70: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/$exit
      -- CP-element group 70: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2762/if_stmt_3220_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2762/if_stmt_3220_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2762/if_stmt_3220_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2762/if_stmt_3220_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2762/R_cmp92_3221_place
      -- CP-element group 70: 	 branch_block_stmt_2762/if_stmt_3220_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2762/if_stmt_3220_else_link/$entry
      -- 
    ca_8767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3213_inst_ack_1, ack => convTransposeD_CP_7773_elements(70)); -- 
    branch_req_8775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(70), ack => if_stmt_3220_branch_req_0); -- 
    -- CP-element group 71:  merge  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2762/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2762/merge_stmt_3226__exit__
      -- CP-element group 71: 	 branch_block_stmt_2762/assign_stmt_3230__entry__
      -- CP-element group 71: 	 branch_block_stmt_2762/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2762/merge_stmt_3226_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2762/merge_stmt_3226_PhiAck/dummy
      -- CP-element group 71: 	 branch_block_stmt_2762/if_stmt_3220_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2762/merge_stmt_3226_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2762/if_stmt_3220_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2762/merge_stmt_3226_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2762/ifx_xend_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2762/assign_stmt_3230/$entry
      -- CP-element group 71: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_Sample/req
      -- 
    if_choice_transition_8780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3220_branch_ack_1, ack => convTransposeD_CP_7773_elements(71)); -- 
    req_8797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(71), ack => WPIPE_Block3_done_3228_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	86 
    -- CP-element group 72: 	82 
    -- CP-element group 72: 	83 
    -- CP-element group 72: 	85 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_2762/if_stmt_3220_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2762/if_stmt_3220_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3220_branch_ack_0, ack => convTransposeD_CP_7773_elements(72)); -- 
    rr_8871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(72), ack => type_cast_2913_inst_req_0); -- 
    cr_8876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(72), ack => type_cast_2913_inst_req_1); -- 
    rr_8894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(72), ack => type_cast_2919_inst_req_0); -- 
    cr_8899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(72), ack => type_cast_2919_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_Update/req
      -- 
    ack_8798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3228_inst_ack_0, ack => convTransposeD_CP_7773_elements(73)); -- 
    req_8802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(73), ack => WPIPE_Block3_done_3228_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2762/$exit
      -- CP-element group 74: 	 branch_block_stmt_2762/branch_block_stmt_2762__exit__
      -- CP-element group 74: 	 branch_block_stmt_2762/assign_stmt_3230__exit__
      -- CP-element group 74: 	 branch_block_stmt_2762/return__
      -- CP-element group 74: 	 branch_block_stmt_2762/merge_stmt_3232__exit__
      -- CP-element group 74: 	 branch_block_stmt_2762/merge_stmt_3232_PhiAck/dummy
      -- CP-element group 74: 	 branch_block_stmt_2762/merge_stmt_3232_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2762/merge_stmt_3232_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2762/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2762/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2762/merge_stmt_3232_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2762/assign_stmt_3230/$exit
      -- CP-element group 74: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2762/assign_stmt_3230/WPIPE_Block3_done_3228_Update/ack
      -- 
    ack_8803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3228_inst_ack_1, ack => convTransposeD_CP_7773_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	33 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Sample/ra
      -- 
    ra_8823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2911_inst_ack_0, ack => convTransposeD_CP_7773_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	33 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Update/ca
      -- 
    ca_8828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2911_inst_ack_1, ack => convTransposeD_CP_7773_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/$exit
      -- CP-element group 77: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/$exit
      -- CP-element group 77: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_req
      -- 
    phi_stmt_2908_req_8829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2908_req_8829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(77), ack => phi_stmt_2908_req_0); -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(75) & convTransposeD_CP_7773_elements(76);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	33 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/ra
      -- 
    ra_8846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2917_inst_ack_0, ack => convTransposeD_CP_7773_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	33 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/ca
      -- 
    ca_8851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2917_inst_ack_1, ack => convTransposeD_CP_7773_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/$exit
      -- CP-element group 80: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/$exit
      -- CP-element group 80: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_req
      -- 
    phi_stmt_2914_req_8852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2914_req_8852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(80), ack => phi_stmt_2914_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(78) & convTransposeD_CP_7773_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	89 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2762/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(77) & convTransposeD_CP_7773_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	72 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Sample/ra
      -- 
    ra_8872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2913_inst_ack_0, ack => convTransposeD_CP_7773_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	72 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Update/ca
      -- 
    ca_8877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2913_inst_ack_1, ack => convTransposeD_CP_7773_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	88 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/$exit
      -- CP-element group 84: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/$exit
      -- CP-element group 84: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2908/phi_stmt_2908_req
      -- 
    phi_stmt_2908_req_8878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2908_req_8878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(84), ack => phi_stmt_2908_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(82) & convTransposeD_CP_7773_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	72 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/ra
      -- 
    ra_8895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2919_inst_ack_0, ack => convTransposeD_CP_7773_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	72 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/ca
      -- 
    ca_8900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2919_inst_ack_1, ack => convTransposeD_CP_7773_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/$exit
      -- CP-element group 87: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/$exit
      -- CP-element group 87: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2914/phi_stmt_2914_req
      -- 
    phi_stmt_2914_req_8901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2914_req_8901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(87), ack => phi_stmt_2914_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(86) & convTransposeD_CP_7773_elements(85);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: 	84 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2762/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(87) & convTransposeD_CP_7773_elements(84);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  merge  fork  transition  place  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	81 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2762/merge_stmt_2907_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_2762/merge_stmt_2907_PhiAck/$entry
      -- 
    convTransposeD_CP_7773_elements(89) <= OrReduce(convTransposeD_CP_7773_elements(81) & convTransposeD_CP_7773_elements(88));
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2762/merge_stmt_2907_PhiAck/phi_stmt_2908_ack
      -- 
    phi_stmt_2908_ack_8906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2908_ack_0, ack => convTransposeD_CP_7773_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_2762/merge_stmt_2907_PhiAck/phi_stmt_2914_ack
      -- 
    phi_stmt_2914_ack_8907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2914_ack_0, ack => convTransposeD_CP_7773_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  place  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	36 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	35 
    -- CP-element group 92: 	34 
    -- CP-element group 92:  members (16) 
      -- CP-element group 92: 	 branch_block_stmt_2762/merge_stmt_2907__exit__
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032__entry__
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/$entry
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2924_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2762/assign_stmt_2925_to_assign_stmt_3032/type_cast_2929_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2762/merge_stmt_2907_PhiAck/$exit
      -- 
    rr_8404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(92), ack => type_cast_2924_inst_req_0); -- 
    cr_8409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(92), ack => type_cast_2924_inst_req_1); -- 
    rr_8418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(92), ack => type_cast_2929_inst_req_0); -- 
    cr_8423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(92), ack => type_cast_2929_inst_req_1); -- 
    convTransposeD_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(90) & convTransposeD_CP_7773_elements(91);
      gj_convTransposeD_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	61 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/Sample/ra
      -- 
    ra_8927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3041_inst_ack_0, ack => convTransposeD_CP_7773_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	61 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/Update/ca
      -- 
    ca_8932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3041_inst_ack_1, ack => convTransposeD_CP_7773_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 95: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/$exit
      -- CP-element group 95: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/$exit
      -- CP-element group 95: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3041/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_2762/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_req
      -- 
    phi_stmt_3035_req_8933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3035_req_8933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(95), ack => phi_stmt_3035_req_1); -- 
    convTransposeD_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(93) & convTransposeD_CP_7773_elements(94);
      gj_convTransposeD_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  output  delay-element  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	38 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 96: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3035/$exit
      -- CP-element group 96: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_sources/type_cast_3039_konst_delay_trans
      -- CP-element group 96: 	 branch_block_stmt_2762/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3035/phi_stmt_3035_req
      -- 
    phi_stmt_3035_req_8944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3035_req_8944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(96), ack => phi_stmt_3035_req_0); -- 
    -- Element group convTransposeD_CP_7773_elements(96) is a control-delay.
    cp_element_96_delay: control_delay_element  generic map(name => " 96_delay", delay_value => 1)  port map(req => convTransposeD_CP_7773_elements(38), ack => convTransposeD_CP_7773_elements(96), clk => clk, reset =>reset);
    -- CP-element group 97:  merge  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_2762/merge_stmt_3034_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_2762/merge_stmt_3034_PhiAck/$entry
      -- 
    convTransposeD_CP_7773_elements(97) <= OrReduce(convTransposeD_CP_7773_elements(95) & convTransposeD_CP_7773_elements(96));
    -- CP-element group 98:  fork  transition  place  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	48 
    -- CP-element group 98: 	57 
    -- CP-element group 98: 	52 
    -- CP-element group 98: 	50 
    -- CP-element group 98: 	44 
    -- CP-element group 98: 	39 
    -- CP-element group 98: 	40 
    -- CP-element group 98: 	59 
    -- CP-element group 98: 	42 
    -- CP-element group 98: 	46 
    -- CP-element group 98: 	54 
    -- CP-element group 98: 	58 
    -- CP-element group 98:  members (45) 
      -- CP-element group 98: 	 branch_block_stmt_2762/merge_stmt_3034__exit__
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140__entry__
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3051_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3081_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3087_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3088_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3092_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3112_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/array_obj_ref_3118_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/addr_of_3119_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/ptr_deref_3122_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2762/assign_stmt_3048_to_assign_stmt_3140/type_cast_3128_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2762/merge_stmt_3034_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_2762/merge_stmt_3034_PhiAck/phi_stmt_3035_ack
      -- 
    phi_stmt_3035_ack_8949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3035_ack_0, ack => convTransposeD_CP_7773_elements(98)); -- 
    rr_8435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => type_cast_3051_inst_req_0); -- 
    cr_8440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => type_cast_3051_inst_req_1); -- 
    cr_8454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => type_cast_3081_inst_req_1); -- 
    req_8485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => array_obj_ref_3087_index_offset_req_1); -- 
    req_8500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => addr_of_3088_final_reg_req_1); -- 
    cr_8545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => ptr_deref_3092_load_0_req_1); -- 
    cr_8564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => type_cast_3112_inst_req_1); -- 
    req_8595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => array_obj_ref_3118_index_offset_req_1); -- 
    req_8610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => addr_of_3119_final_reg_req_1); -- 
    cr_8660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => ptr_deref_3122_store_0_req_1); -- 
    rr_8669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => type_cast_3128_inst_req_0); -- 
    cr_8674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(98), ack => type_cast_3128_inst_req_1); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	66 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/Sample/ra
      -- 
    ra_9001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3206_inst_ack_0, ack => convTransposeD_CP_7773_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	66 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/Update/ca
      -- 
    ca_9006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3206_inst_ack_1, ack => convTransposeD_CP_7773_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	105 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/$exit
      -- CP-element group 101: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/$exit
      -- CP-element group 101: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3206/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_req
      -- 
    phi_stmt_3203_req_9007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3203_req_9007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(101), ack => phi_stmt_3203_req_0); -- 
    convTransposeD_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(99) & convTransposeD_CP_7773_elements(100);
      gj_convTransposeD_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/Sample/ra
      -- 
    ra_9024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3200_inst_ack_0, ack => convTransposeD_CP_7773_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/Update/ca
      -- 
    ca_9029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3200_inst_ack_1, ack => convTransposeD_CP_7773_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/$exit
      -- CP-element group 104: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/$exit
      -- CP-element group 104: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3200/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_req
      -- 
    phi_stmt_3197_req_9030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3197_req_9030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(104), ack => phi_stmt_3197_req_0); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(102) & convTransposeD_CP_7773_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	101 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	113 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2762/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(101) & convTransposeD_CP_7773_elements(104);
      gj_convTransposeD_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	68 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/Sample/ra
      -- 
    ra_9050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3208_inst_ack_0, ack => convTransposeD_CP_7773_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	68 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/Update/ca
      -- 
    ca_9055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3208_inst_ack_1, ack => convTransposeD_CP_7773_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/$exit
      -- CP-element group 108: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/$exit
      -- CP-element group 108: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_sources/type_cast_3208/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3203/phi_stmt_3203_req
      -- 
    phi_stmt_3203_req_9056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3203_req_9056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(108), ack => phi_stmt_3203_req_1); -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(106) & convTransposeD_CP_7773_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	68 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/Sample/ra
      -- 
    ra_9073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3202_inst_ack_0, ack => convTransposeD_CP_7773_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	68 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/Update/ca
      -- 
    ca_9078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3202_inst_ack_1, ack => convTransposeD_CP_7773_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/$exit
      -- CP-element group 111: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/$exit
      -- CP-element group 111: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_sources/type_cast_3202/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3197/phi_stmt_3197_req
      -- 
    phi_stmt_3197_req_9079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3197_req_9079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(111), ack => phi_stmt_3197_req_1); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(109) & convTransposeD_CP_7773_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2762/ifx_xthen83_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(108) & convTransposeD_CP_7773_elements(111);
      gj_convTransposeD_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  merge  fork  transition  place  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	105 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2762/merge_stmt_3196_PhiReqMerge
      -- CP-element group 113: 	 branch_block_stmt_2762/merge_stmt_3196_PhiAck/$entry
      -- 
    convTransposeD_CP_7773_elements(113) <= OrReduce(convTransposeD_CP_7773_elements(105) & convTransposeD_CP_7773_elements(112));
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2762/merge_stmt_3196_PhiAck/phi_stmt_3197_ack
      -- 
    phi_stmt_3197_ack_9084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3197_ack_0, ack => convTransposeD_CP_7773_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2762/merge_stmt_3196_PhiAck/phi_stmt_3203_ack
      -- 
    phi_stmt_3203_ack_9085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3203_ack_0, ack => convTransposeD_CP_7773_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: 	70 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_2762/merge_stmt_3196__exit__
      -- CP-element group 116: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219__entry__
      -- CP-element group 116: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/$entry
      -- CP-element group 116: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_update_start_
      -- CP-element group 116: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_2762/assign_stmt_3214_to_assign_stmt_3219/type_cast_3213_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_2762/merge_stmt_3196_PhiAck/$exit
      -- 
    rr_8761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(116), ack => type_cast_3213_inst_req_0); -- 
    cr_8766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7773_elements(116), ack => type_cast_3213_inst_req_1); -- 
    convTransposeD_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7773_elements(114) & convTransposeD_CP_7773_elements(115);
      gj_convTransposeD_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7773_elements(116), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2994_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3015_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3075_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3106_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2850_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2850_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom65_3117_resized : std_logic_vector(13 downto 0);
    signal R_idxprom65_3117_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3086_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3086_scaled : std_logic_vector(13 downto 0);
    signal add21_3057 : std_logic_vector(31 downto 0);
    signal add29_2955 : std_logic_vector(31 downto 0);
    signal add40_2970 : std_logic_vector(31 downto 0);
    signal add55_3027 : std_logic_vector(31 downto 0);
    signal add57_3062 : std_logic_vector(31 downto 0);
    signal add70_3135 : std_logic_vector(31 downto 0);
    signal add_2940 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3087_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3087_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3087_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3087_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3087_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3087_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3118_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3118_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3118_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3118_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3118_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3118_root_address : std_logic_vector(13 downto 0);
    signal arrayidx66_3120 : std_logic_vector(31 downto 0);
    signal arrayidx_3089 : std_logic_vector(31 downto 0);
    signal call_2765 : std_logic_vector(15 downto 0);
    signal cmp81_3171 : std_logic_vector(0 downto 0);
    signal cmp92_3219 : std_logic_vector(0 downto 0);
    signal cmp_3140 : std_logic_vector(0 downto 0);
    signal conv13105_3052 : std_logic_vector(31 downto 0);
    signal conv16_2925 : std_logic_vector(31 downto 0);
    signal conv19_2930 : std_logic_vector(31 downto 0);
    signal conv26_2836 : std_logic_vector(31 downto 0);
    signal conv31_2855 : std_logic_vector(31 downto 0);
    signal conv37_2869 : std_logic_vector(31 downto 0);
    signal conv4_2810 : std_logic_vector(15 downto 0);
    signal conv50_2996 : std_logic_vector(31 downto 0);
    signal conv53_3017 : std_logic_vector(31 downto 0);
    signal conv69_3129 : std_logic_vector(31 downto 0);
    signal conv79_3166 : std_logic_vector(31 downto 0);
    signal conv88_3194 : std_logic_vector(15 downto 0);
    signal conv90_3214 : std_logic_vector(31 downto 0);
    signal conv_2788 : std_logic_vector(15 downto 0);
    signal div3_2806 : std_logic_vector(31 downto 0);
    signal div87_3190 : std_logic_vector(31 downto 0);
    signal div_2784 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2901 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2774 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2796 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2818 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2828 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2844 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2861 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2877 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2889 : std_logic_vector(31 downto 0);
    signal idxprom65_3113 : std_logic_vector(63 downto 0);
    signal idxprom_3082 : std_logic_vector(63 downto 0);
    signal inc85_3184 : std_logic_vector(15 downto 0);
    signal inc_3161 : std_logic_vector(15 downto 0);
    signal indvar_3035 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_3153 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_3203 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2914 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2908 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_3197 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_3048 : std_logic_vector(15 downto 0);
    signal mul20_2945 : std_logic_vector(31 downto 0);
    signal mul27_2950 : std_logic_vector(31 downto 0);
    signal mul38_2965 : std_logic_vector(31 downto 0);
    signal mul54_3022 : std_logic_vector(31 downto 0);
    signal mul56_3032 : std_logic_vector(31 downto 0);
    signal mul_2935 : std_logic_vector(31 downto 0);
    signal ptr_deref_2777_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2777_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2777_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2777_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2777_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2799_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2799_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2799_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2799_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2799_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2821_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2821_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2821_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2821_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2821_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2831_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2831_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2831_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2831_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2831_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2847_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2847_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2847_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2847_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2847_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2864_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2864_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2864_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2864_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2864_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2880_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2880_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2880_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2880_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2880_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2892_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2892_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2892_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2892_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2892_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2904_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2904_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2904_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2904_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2904_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3092_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3092_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3092_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3092_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3092_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3122_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3122_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3122_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3122_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3122_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3122_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext106_3008 : std_logic_vector(31 downto 0);
    signal sext108_3068 : std_logic_vector(31 downto 0);
    signal sext109_3099 : std_logic_vector(31 downto 0);
    signal sext_2987 : std_logic_vector(31 downto 0);
    signal shr64_3108 : std_logic_vector(31 downto 0);
    signal shr_3077 : std_logic_vector(31 downto 0);
    signal sub32_3002 : std_logic_vector(31 downto 0);
    signal sub43_2975 : std_logic_vector(31 downto 0);
    signal sub44_2981 : std_logic_vector(31 downto 0);
    signal sub_2960 : std_logic_vector(31 downto 0);
    signal tmp14_2822 : std_logic_vector(31 downto 0);
    signal tmp25_2832 : std_logic_vector(15 downto 0);
    signal tmp28_2848 : std_logic_vector(31 downto 0);
    signal tmp2_2800 : std_logic_vector(31 downto 0);
    signal tmp30_2851 : std_logic_vector(15 downto 0);
    signal tmp36_2865 : std_logic_vector(15 downto 0);
    signal tmp39_2881 : std_logic_vector(31 downto 0);
    signal tmp48_2893 : std_logic_vector(31 downto 0);
    signal tmp51_2905 : std_logic_vector(31 downto 0);
    signal tmp61_3093 : std_logic_vector(63 downto 0);
    signal tmp_2778 : std_logic_vector(31 downto 0);
    signal type_cast_2782_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2804_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2911_wire : std_logic_vector(15 downto 0);
    signal type_cast_2913_wire : std_logic_vector(15 downto 0);
    signal type_cast_2917_wire : std_logic_vector(15 downto 0);
    signal type_cast_2919_wire : std_logic_vector(15 downto 0);
    signal type_cast_2923_wire : std_logic_vector(31 downto 0);
    signal type_cast_2928_wire : std_logic_vector(31 downto 0);
    signal type_cast_2979_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2985_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2990_wire : std_logic_vector(31 downto 0);
    signal type_cast_2993_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3000_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3006_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3011_wire : std_logic_vector(31 downto 0);
    signal type_cast_3014_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3039_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3041_wire : std_logic_vector(15 downto 0);
    signal type_cast_3046_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3066_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3071_wire : std_logic_vector(31 downto 0);
    signal type_cast_3074_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3080_wire : std_logic_vector(63 downto 0);
    signal type_cast_3097_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3102_wire : std_logic_vector(31 downto 0);
    signal type_cast_3105_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3111_wire : std_logic_vector(63 downto 0);
    signal type_cast_3127_wire : std_logic_vector(31 downto 0);
    signal type_cast_3133_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3151_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3159_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3164_wire : std_logic_vector(31 downto 0);
    signal type_cast_3182_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3188_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3200_wire : std_logic_vector(15 downto 0);
    signal type_cast_3202_wire : std_logic_vector(15 downto 0);
    signal type_cast_3206_wire : std_logic_vector(15 downto 0);
    signal type_cast_3208_wire : std_logic_vector(15 downto 0);
    signal type_cast_3212_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2850_word_address_0 <= "0";
    array_obj_ref_3087_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3087_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3087_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3087_resized_base_address <= "00000000000000";
    array_obj_ref_3118_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3118_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3118_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3118_resized_base_address <= "00000000000000";
    iNsTr_10_2901 <= "00000000000000000000000000000011";
    iNsTr_2_2774 <= "00000000000000000000000000000010";
    iNsTr_3_2796 <= "00000000000000000000000000000011";
    iNsTr_4_2818 <= "00000000000000000000000000000100";
    iNsTr_5_2828 <= "00000000000000000000000000000000";
    iNsTr_6_2844 <= "00000000000000000000000000000011";
    iNsTr_7_2861 <= "00000000000000000000000000000001";
    iNsTr_8_2877 <= "00000000000000000000000000000100";
    iNsTr_9_2889 <= "00000000000000000000000000000100";
    ptr_deref_2777_word_offset_0 <= "0000000";
    ptr_deref_2799_word_offset_0 <= "0000000";
    ptr_deref_2821_word_offset_0 <= "0000000";
    ptr_deref_2831_word_offset_0 <= "0";
    ptr_deref_2847_word_offset_0 <= "0000000";
    ptr_deref_2864_word_offset_0 <= "0";
    ptr_deref_2880_word_offset_0 <= "0000000";
    ptr_deref_2892_word_offset_0 <= "0000000";
    ptr_deref_2904_word_offset_0 <= "0000000";
    ptr_deref_3092_word_offset_0 <= "00000000000000";
    ptr_deref_3122_word_offset_0 <= "00000000000000";
    type_cast_2782_wire_constant <= "00000000000000000000000000000001";
    type_cast_2804_wire_constant <= "00000000000000000000000000000001";
    type_cast_2979_wire_constant <= "00000000000000000000000000010000";
    type_cast_2985_wire_constant <= "11111111111111110000000000000000";
    type_cast_2993_wire_constant <= "00000000000000000000000000010000";
    type_cast_3000_wire_constant <= "00000000000000000000000000010000";
    type_cast_3006_wire_constant <= "11111111111111110000000000000000";
    type_cast_3014_wire_constant <= "00000000000000000000000000010000";
    type_cast_3039_wire_constant <= "0000000000000000";
    type_cast_3046_wire_constant <= "0000000000000100";
    type_cast_3066_wire_constant <= "00000000000000000000000000010000";
    type_cast_3074_wire_constant <= "00000000000000000000000000010010";
    type_cast_3097_wire_constant <= "00000000000000000000000000010000";
    type_cast_3105_wire_constant <= "00000000000000000000000000010010";
    type_cast_3133_wire_constant <= "00000000000000000000000000000100";
    type_cast_3151_wire_constant <= "0000000000000001";
    type_cast_3159_wire_constant <= "0000000000000001";
    type_cast_3182_wire_constant <= "0000000000000001";
    type_cast_3188_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_2908: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2911_wire & type_cast_2913_wire;
      req <= phi_stmt_2908_req_0 & phi_stmt_2908_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2908",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2908_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2908,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2908
    phi_stmt_2914: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2917_wire & type_cast_2919_wire;
      req <= phi_stmt_2914_req_0 & phi_stmt_2914_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2914",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2914_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2914,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2914
    phi_stmt_3035: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3039_wire_constant & type_cast_3041_wire;
      req <= phi_stmt_3035_req_0 & phi_stmt_3035_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3035",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3035_ack_0,
          idata => idata,
          odata => indvar_3035,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3035
    phi_stmt_3197: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3200_wire & type_cast_3202_wire;
      req <= phi_stmt_3197_req_0 & phi_stmt_3197_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3197",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3197_ack_0,
          idata => idata,
          odata => input_dim1x_x2_3197,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3197
    phi_stmt_3203: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3206_wire & type_cast_3208_wire;
      req <= phi_stmt_3203_req_0 & phi_stmt_3203_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3203",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3203_ack_0,
          idata => idata,
          odata => input_dim0x_x0_3203,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3203
    addr_of_3088_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3088_final_reg_req_0;
      addr_of_3088_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3088_final_reg_req_1;
      addr_of_3088_final_reg_ack_1<= rack(0);
      addr_of_3088_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3088_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3087_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_3089,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3119_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3119_final_reg_req_0;
      addr_of_3119_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3119_final_reg_req_1;
      addr_of_3119_final_reg_ack_1<= rack(0);
      addr_of_3119_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3119_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3118_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx66_3120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2787_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2787_inst_req_0;
      type_cast_2787_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2787_inst_req_1;
      type_cast_2787_inst_ack_1<= rack(0);
      type_cast_2787_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2787_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2784,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2809_inst_req_0;
      type_cast_2809_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2809_inst_req_1;
      type_cast_2809_inst_ack_1<= rack(0);
      type_cast_2809_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div3_2806,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_2810,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2835_inst_req_0;
      type_cast_2835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2835_inst_req_1;
      type_cast_2835_inst_ack_1<= rack(0);
      type_cast_2835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp25_2832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_2836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2854_inst_req_0;
      type_cast_2854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2854_inst_req_1;
      type_cast_2854_inst_ack_1<= rack(0);
      type_cast_2854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp30_2851,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_2855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2868_inst_req_0;
      type_cast_2868_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2868_inst_req_1;
      type_cast_2868_inst_ack_1<= rack(0);
      type_cast_2868_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2868_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp36_2865,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_2869,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2911_inst_req_0;
      type_cast_2911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2911_inst_req_1;
      type_cast_2911_inst_ack_1<= rack(0);
      type_cast_2911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2911_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_2810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2911_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2913_inst_req_0;
      type_cast_2913_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2913_inst_req_1;
      type_cast_2913_inst_ack_1<= rack(0);
      type_cast_2913_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2913_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_3197,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2913_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2917_inst_req_0;
      type_cast_2917_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2917_inst_req_1;
      type_cast_2917_inst_ack_1<= rack(0);
      type_cast_2917_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2788,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2917_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2919_inst_req_0;
      type_cast_2919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2919_inst_req_1;
      type_cast_2919_inst_ack_1<= rack(0);
      type_cast_2919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_3203,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2919_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2924_inst_req_0;
      type_cast_2924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2924_inst_req_1;
      type_cast_2924_inst_ack_1<= rack(0);
      type_cast_2924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2923_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2929_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2929_inst_req_0;
      type_cast_2929_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2929_inst_req_1;
      type_cast_2929_inst_ack_1<= rack(0);
      type_cast_2929_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2929_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2928_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_2930,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2990_inst
    process(sext_2987) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2987(31 downto 0);
      type_cast_2990_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2995_inst
    process(ASHR_i32_i32_2994_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2994_wire(31 downto 0);
      conv50_2996 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3011_inst
    process(sext106_3008) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_3008(31 downto 0);
      type_cast_3011_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3016_inst
    process(ASHR_i32_i32_3015_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3015_wire(31 downto 0);
      conv53_3017 <= tmp_var; -- 
    end process;
    type_cast_3041_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3041_inst_req_0;
      type_cast_3041_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3041_inst_req_1;
      type_cast_3041_inst_ack_1<= rack(0);
      type_cast_3041_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3041_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_3153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3041_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3051_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3051_inst_req_0;
      type_cast_3051_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3051_inst_req_1;
      type_cast_3051_inst_ack_1<= rack(0);
      type_cast_3051_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3051_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_3048,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13105_3052,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3071_inst
    process(sext108_3068) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext108_3068(31 downto 0);
      type_cast_3071_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3076_inst
    process(ASHR_i32_i32_3075_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3075_wire(31 downto 0);
      shr_3077 <= tmp_var; -- 
    end process;
    type_cast_3081_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3081_inst_req_0;
      type_cast_3081_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3081_inst_req_1;
      type_cast_3081_inst_ack_1<= rack(0);
      type_cast_3081_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3081_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3080_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3082,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3102_inst
    process(sext109_3099) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext109_3099(31 downto 0);
      type_cast_3102_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3107_inst
    process(ASHR_i32_i32_3106_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3106_wire(31 downto 0);
      shr64_3108 <= tmp_var; -- 
    end process;
    type_cast_3112_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3112_inst_req_0;
      type_cast_3112_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3112_inst_req_1;
      type_cast_3112_inst_ack_1<= rack(0);
      type_cast_3112_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3112_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3111_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom65_3113,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3128_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3128_inst_req_0;
      type_cast_3128_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3128_inst_req_1;
      type_cast_3128_inst_ack_1<= rack(0);
      type_cast_3128_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3128_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3127_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_3129,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3165_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3165_inst_req_0;
      type_cast_3165_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3165_inst_req_1;
      type_cast_3165_inst_ack_1<= rack(0);
      type_cast_3165_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3165_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3164_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_3166,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3193_inst_req_0;
      type_cast_3193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3193_inst_req_1;
      type_cast_3193_inst_ack_1<= rack(0);
      type_cast_3193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div87_3190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_3194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3200_inst_req_0;
      type_cast_3200_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3200_inst_req_1;
      type_cast_3200_inst_ack_1<= rack(0);
      type_cast_3200_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3200_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_3161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3200_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3202_inst_req_0;
      type_cast_3202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3202_inst_req_1;
      type_cast_3202_inst_ack_1<= rack(0);
      type_cast_3202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv88_3194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3202_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3206_inst_req_0;
      type_cast_3206_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3206_inst_req_1;
      type_cast_3206_inst_ack_1<= rack(0);
      type_cast_3206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_2914,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3206_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3208_inst_req_0;
      type_cast_3208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3208_inst_req_1;
      type_cast_3208_inst_ack_1<= rack(0);
      type_cast_3208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc85_3184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3208_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3213_inst_req_0;
      type_cast_3213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3213_inst_req_1;
      type_cast_3213_inst_ack_1<= rack(0);
      type_cast_3213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3212_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_3214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2850_gather_scatter
    process(LOAD_padding_2850_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2850_data_0;
      ov(15 downto 0) := iv;
      tmp30_2851 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3087_index_1_rename
    process(R_idxprom_3086_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3086_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3086_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3087_index_1_resize
    process(idxprom_3082) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3082;
      ov := iv(13 downto 0);
      R_idxprom_3086_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3087_root_address_inst
    process(array_obj_ref_3087_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3087_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3087_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3118_index_1_rename
    process(R_idxprom65_3117_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom65_3117_resized;
      ov(13 downto 0) := iv;
      R_idxprom65_3117_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3118_index_1_resize
    process(idxprom65_3113) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom65_3113;
      ov := iv(13 downto 0);
      R_idxprom65_3117_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3118_root_address_inst
    process(array_obj_ref_3118_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3118_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3118_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2777_addr_0
    process(ptr_deref_2777_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2777_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2777_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2777_base_resize
    process(iNsTr_2_2774) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2774;
      ov := iv(6 downto 0);
      ptr_deref_2777_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2777_gather_scatter
    process(ptr_deref_2777_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2777_data_0;
      ov(31 downto 0) := iv;
      tmp_2778 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2777_root_address_inst
    process(ptr_deref_2777_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2777_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2777_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2799_addr_0
    process(ptr_deref_2799_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2799_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2799_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2799_base_resize
    process(iNsTr_3_2796) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2796;
      ov := iv(6 downto 0);
      ptr_deref_2799_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2799_gather_scatter
    process(ptr_deref_2799_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2799_data_0;
      ov(31 downto 0) := iv;
      tmp2_2800 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2799_root_address_inst
    process(ptr_deref_2799_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2799_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2799_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2821_addr_0
    process(ptr_deref_2821_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2821_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2821_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2821_base_resize
    process(iNsTr_4_2818) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2818;
      ov := iv(6 downto 0);
      ptr_deref_2821_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2821_gather_scatter
    process(ptr_deref_2821_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2821_data_0;
      ov(31 downto 0) := iv;
      tmp14_2822 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2821_root_address_inst
    process(ptr_deref_2821_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2821_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2821_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2831_addr_0
    process(ptr_deref_2831_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2831_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2831_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2831_base_resize
    process(iNsTr_5_2828) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2828;
      ov := iv(0 downto 0);
      ptr_deref_2831_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2831_gather_scatter
    process(ptr_deref_2831_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2831_data_0;
      ov(15 downto 0) := iv;
      tmp25_2832 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2831_root_address_inst
    process(ptr_deref_2831_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2831_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2831_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2847_addr_0
    process(ptr_deref_2847_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2847_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2847_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2847_base_resize
    process(iNsTr_6_2844) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2844;
      ov := iv(6 downto 0);
      ptr_deref_2847_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2847_gather_scatter
    process(ptr_deref_2847_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2847_data_0;
      ov(31 downto 0) := iv;
      tmp28_2848 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2847_root_address_inst
    process(ptr_deref_2847_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2847_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2847_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2864_addr_0
    process(ptr_deref_2864_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2864_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2864_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2864_base_resize
    process(iNsTr_7_2861) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2861;
      ov := iv(0 downto 0);
      ptr_deref_2864_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2864_gather_scatter
    process(ptr_deref_2864_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2864_data_0;
      ov(15 downto 0) := iv;
      tmp36_2865 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2864_root_address_inst
    process(ptr_deref_2864_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2864_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2864_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2880_addr_0
    process(ptr_deref_2880_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2880_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2880_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2880_base_resize
    process(iNsTr_8_2877) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2877;
      ov := iv(6 downto 0);
      ptr_deref_2880_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2880_gather_scatter
    process(ptr_deref_2880_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2880_data_0;
      ov(31 downto 0) := iv;
      tmp39_2881 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2880_root_address_inst
    process(ptr_deref_2880_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2880_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2880_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2892_addr_0
    process(ptr_deref_2892_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2892_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2892_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2892_base_resize
    process(iNsTr_9_2889) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2889;
      ov := iv(6 downto 0);
      ptr_deref_2892_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2892_gather_scatter
    process(ptr_deref_2892_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2892_data_0;
      ov(31 downto 0) := iv;
      tmp48_2893 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2892_root_address_inst
    process(ptr_deref_2892_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2892_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2892_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2904_addr_0
    process(ptr_deref_2904_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2904_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2904_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2904_base_resize
    process(iNsTr_10_2901) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2901;
      ov := iv(6 downto 0);
      ptr_deref_2904_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2904_gather_scatter
    process(ptr_deref_2904_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2904_data_0;
      ov(31 downto 0) := iv;
      tmp51_2905 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2904_root_address_inst
    process(ptr_deref_2904_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2904_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2904_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3092_addr_0
    process(ptr_deref_3092_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3092_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3092_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3092_base_resize
    process(arrayidx_3089) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_3089;
      ov := iv(13 downto 0);
      ptr_deref_3092_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3092_gather_scatter
    process(ptr_deref_3092_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3092_data_0;
      ov(63 downto 0) := iv;
      tmp61_3093 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3092_root_address_inst
    process(ptr_deref_3092_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3092_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3092_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3122_addr_0
    process(ptr_deref_3122_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3122_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3122_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3122_base_resize
    process(arrayidx66_3120) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx66_3120;
      ov := iv(13 downto 0);
      ptr_deref_3122_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3122_gather_scatter
    process(tmp61_3093) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp61_3093;
      ov(63 downto 0) := iv;
      ptr_deref_3122_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3122_root_address_inst
    process(ptr_deref_3122_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3122_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3122_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3141_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_3140;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3141_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3141_branch_req_0,
          ack0 => if_stmt_3141_branch_ack_0,
          ack1 => if_stmt_3141_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3172_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp81_3171;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3172_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3172_branch_req_0,
          ack0 => if_stmt_3172_branch_ack_0,
          ack1 => if_stmt_3172_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3220_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp92_3219;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3220_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3220_branch_req_0,
          ack0 => if_stmt_3220_branch_ack_0,
          ack1 => if_stmt_3220_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3152_inst
    process(indvar_3035) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_3035, type_cast_3151_wire_constant, tmp_var);
      indvarx_xnext_3153 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3160_inst
    process(input_dim1x_x1x_xph_2908) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2908, type_cast_3159_wire_constant, tmp_var);
      inc_3161 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3183_inst
    process(input_dim0x_x2x_xph_2914) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_2914, type_cast_3182_wire_constant, tmp_var);
      inc85_3184 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2939_inst
    process(mul_2935, conv16_2925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2935, conv16_2925, tmp_var);
      add_2940 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2954_inst
    process(mul27_2950, tmp28_2848) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul27_2950, tmp28_2848, tmp_var);
      add29_2955 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2969_inst
    process(mul38_2965, tmp39_2881) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul38_2965, tmp39_2881, tmp_var);
      add40_2970 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2986_inst
    process(sub44_2981) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub44_2981, type_cast_2985_wire_constant, tmp_var);
      sext_2987 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3007_inst
    process(sub32_3002) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub32_3002, type_cast_3006_wire_constant, tmp_var);
      sext106_3008 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3026_inst
    process(conv50_2996, mul54_3022) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv50_2996, mul54_3022, tmp_var);
      add55_3027 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3056_inst
    process(mul20_2945, conv13105_3052) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul20_2945, conv13105_3052, tmp_var);
      add21_3057 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3061_inst
    process(mul56_3032, conv13105_3052) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul56_3032, conv13105_3052, tmp_var);
      add57_3062 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3134_inst
    process(conv69_3129) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv69_3129, type_cast_3133_wire_constant, tmp_var);
      add70_3135 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2994_inst
    process(type_cast_2990_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2990_wire, type_cast_2993_wire_constant, tmp_var);
      ASHR_i32_i32_2994_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3015_inst
    process(type_cast_3011_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3011_wire, type_cast_3014_wire_constant, tmp_var);
      ASHR_i32_i32_3015_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3075_inst
    process(type_cast_3071_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3071_wire, type_cast_3074_wire_constant, tmp_var);
      ASHR_i32_i32_3075_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3106_inst
    process(type_cast_3102_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3102_wire, type_cast_3105_wire_constant, tmp_var);
      ASHR_i32_i32_3106_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3170_inst
    process(conv79_3166, tmp2_2800) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv79_3166, tmp2_2800, tmp_var);
      cmp81_3171 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3218_inst
    process(conv90_3214, tmp_2778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv90_3214, tmp_2778, tmp_var);
      cmp92_3219 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2783_inst
    process(tmp_2778) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2778, type_cast_2782_wire_constant, tmp_var);
      div_2784 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2805_inst
    process(tmp2_2800) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2800, type_cast_2804_wire_constant, tmp_var);
      div3_2806 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3189_inst
    process(tmp2_2800) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2800, type_cast_3188_wire_constant, tmp_var);
      div87_3190 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3047_inst
    process(indvar_3035) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_3035, type_cast_3046_wire_constant, tmp_var);
      input_dim2x_x1_3048 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2934_inst
    process(tmp2_2800, conv19_2930) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_2800, conv19_2930, tmp_var);
      mul_2935 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2944_inst
    process(add_2940, tmp14_2822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2940, tmp14_2822, tmp_var);
      mul20_2945 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2949_inst
    process(conv26_2836, conv19_2930) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv26_2836, conv19_2930, tmp_var);
      mul27_2950 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2964_inst
    process(conv37_2869, conv16_2925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv37_2869, conv16_2925, tmp_var);
      mul38_2965 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3021_inst
    process(tmp51_2905, conv53_3017) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp51_2905, conv53_3017, tmp_var);
      mul54_3022 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3031_inst
    process(add55_3027, tmp48_2893) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add55_3027, tmp48_2893, tmp_var);
      mul56_3032 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2980_inst
    process(sub43_2975) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub43_2975, type_cast_2979_wire_constant, tmp_var);
      sub44_2981 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3001_inst
    process(sub_2960) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2960, type_cast_3000_wire_constant, tmp_var);
      sub32_3002 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3067_inst
    process(add21_3057) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add21_3057, type_cast_3066_wire_constant, tmp_var);
      sext108_3068 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3098_inst
    process(add57_3062) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add57_3062, type_cast_3097_wire_constant, tmp_var);
      sext109_3099 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2959_inst
    process(add29_2955, conv31_2855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add29_2955, conv31_2855, tmp_var);
      sub_2960 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2974_inst
    process(add40_2970, conv31_2855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add40_2970, conv31_2855, tmp_var);
      sub43_2975 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_3139_inst
    process(add70_3135, tmp14_2822) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add70_3135, tmp14_2822, tmp_var);
      cmp_3140 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_3087_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3086_scaled;
      array_obj_ref_3087_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3087_index_offset_req_0;
      array_obj_ref_3087_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3087_index_offset_req_1;
      array_obj_ref_3087_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_3118_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom65_3117_scaled;
      array_obj_ref_3118_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3118_index_offset_req_0;
      array_obj_ref_3118_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3118_index_offset_req_1;
      array_obj_ref_3118_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_2923_inst
    process(input_dim1x_x1x_xph_2908) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2908, tmp_var);
      type_cast_2923_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2928_inst
    process(input_dim0x_x2x_xph_2914) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2914, tmp_var);
      type_cast_2928_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3080_inst
    process(shr_3077) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_3077, tmp_var);
      type_cast_3080_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3111_inst
    process(shr64_3108) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr64_3108, tmp_var);
      type_cast_3111_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3127_inst
    process(input_dim2x_x1_3048) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_3048, tmp_var);
      type_cast_3127_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3164_inst
    process(inc_3161) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3161, tmp_var);
      type_cast_3164_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3212_inst
    process(input_dim0x_x0_3203) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_3203, tmp_var);
      type_cast_3212_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2850_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2850_load_0_req_0;
      LOAD_padding_2850_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2850_load_0_req_1;
      LOAD_padding_2850_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2850_word_address_0;
      LOAD_padding_2850_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2821_load_0 ptr_deref_2777_load_0 ptr_deref_2799_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2821_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2777_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2799_load_0_req_0;
      ptr_deref_2821_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2777_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2799_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2821_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2777_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2799_load_0_req_1;
      ptr_deref_2821_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2777_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2799_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2821_word_address_0 & ptr_deref_2777_word_address_0 & ptr_deref_2799_word_address_0;
      ptr_deref_2821_data_0 <= data_out(95 downto 64);
      ptr_deref_2777_data_0 <= data_out(63 downto 32);
      ptr_deref_2799_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2864_load_0 ptr_deref_2831_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2864_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2831_load_0_req_0;
      ptr_deref_2864_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2831_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2864_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2831_load_0_req_1;
      ptr_deref_2864_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2831_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2864_word_address_0 & ptr_deref_2831_word_address_0;
      ptr_deref_2864_data_0 <= data_out(31 downto 16);
      ptr_deref_2831_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2847_load_0 ptr_deref_2880_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2847_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2880_load_0_req_0;
      ptr_deref_2847_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2880_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2847_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2880_load_0_req_1;
      ptr_deref_2847_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2880_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2847_word_address_0 & ptr_deref_2880_word_address_0;
      ptr_deref_2847_data_0 <= data_out(63 downto 32);
      ptr_deref_2880_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2892_load_0 ptr_deref_2904_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2892_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2904_load_0_req_0;
      ptr_deref_2892_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2904_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2892_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2904_load_0_req_1;
      ptr_deref_2892_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2904_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2892_word_address_0 & ptr_deref_2904_word_address_0;
      ptr_deref_2892_data_0 <= data_out(63 downto 32);
      ptr_deref_2904_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_3092_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3092_load_0_req_0;
      ptr_deref_3092_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3092_load_0_req_1;
      ptr_deref_3092_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3092_word_address_0;
      ptr_deref_3092_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_3122_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3122_store_0_req_0;
      ptr_deref_3122_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3122_store_0_req_1;
      ptr_deref_3122_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3122_word_address_0;
      data_in <= ptr_deref_3122_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2764_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_start_2764_inst_req_0;
      RPIPE_Block3_start_2764_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_start_2764_inst_req_1;
      RPIPE_Block3_start_2764_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2765 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_3228_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_3228_inst_req_0;
      WPIPE_Block3_done_3228_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_3228_inst_req_1;
      WPIPE_Block3_done_3228_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2765;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_3305_start: Boolean;
  signal sendOutput_CP_3305_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1178_inst_req_0 : boolean;
  signal type_cast_1178_inst_ack_0 : boolean;
  signal ptr_deref_1133_load_0_req_1 : boolean;
  signal if_stmt_1151_branch_req_0 : boolean;
  signal ptr_deref_1121_load_0_ack_1 : boolean;
  signal ptr_deref_1212_load_0_ack_0 : boolean;
  signal ptr_deref_1109_load_0_ack_1 : boolean;
  signal array_obj_ref_1207_index_offset_ack_1 : boolean;
  signal ptr_deref_1109_load_0_req_1 : boolean;
  signal ptr_deref_1212_load_0_req_0 : boolean;
  signal ptr_deref_1133_load_0_ack_0 : boolean;
  signal array_obj_ref_1207_index_offset_req_1 : boolean;
  signal ptr_deref_1133_load_0_req_0 : boolean;
  signal addr_of_1208_final_reg_ack_1 : boolean;
  signal type_cast_1178_inst_req_1 : boolean;
  signal type_cast_1246_inst_req_1 : boolean;
  signal type_cast_1216_inst_req_1 : boolean;
  signal type_cast_1216_inst_ack_1 : boolean;
  signal ptr_deref_1133_load_0_ack_1 : boolean;
  signal addr_of_1208_final_reg_req_1 : boolean;
  signal type_cast_1178_inst_ack_1 : boolean;
  signal ptr_deref_1212_load_0_ack_1 : boolean;
  signal type_cast_1216_inst_req_0 : boolean;
  signal type_cast_1216_inst_ack_0 : boolean;
  signal ptr_deref_1121_load_0_req_0 : boolean;
  signal type_cast_1226_inst_req_1 : boolean;
  signal type_cast_1226_inst_ack_1 : boolean;
  signal ptr_deref_1212_load_0_req_1 : boolean;
  signal array_obj_ref_1207_index_offset_ack_0 : boolean;
  signal type_cast_1246_inst_ack_1 : boolean;
  signal ptr_deref_1121_load_0_ack_0 : boolean;
  signal array_obj_ref_1207_index_offset_req_0 : boolean;
  signal ptr_deref_1109_load_0_req_0 : boolean;
  signal type_cast_1246_inst_req_0 : boolean;
  signal type_cast_1246_inst_ack_0 : boolean;
  signal addr_of_1208_final_reg_req_0 : boolean;
  signal type_cast_1226_inst_ack_0 : boolean;
  signal ptr_deref_1109_load_0_ack_0 : boolean;
  signal addr_of_1208_final_reg_ack_0 : boolean;
  signal type_cast_1236_inst_req_1 : boolean;
  signal type_cast_1236_inst_ack_1 : boolean;
  signal if_stmt_1151_branch_ack_1 : boolean;
  signal type_cast_1256_inst_req_0 : boolean;
  signal ptr_deref_1121_load_0_req_1 : boolean;
  signal type_cast_1256_inst_ack_0 : boolean;
  signal type_cast_1256_inst_req_1 : boolean;
  signal type_cast_1256_inst_ack_1 : boolean;
  signal type_cast_1236_inst_ack_0 : boolean;
  signal type_cast_1236_inst_req_0 : boolean;
  signal if_stmt_1151_branch_ack_0 : boolean;
  signal type_cast_1226_inst_req_0 : boolean;
  signal type_cast_1266_inst_req_0 : boolean;
  signal type_cast_1266_inst_ack_0 : boolean;
  signal type_cast_1266_inst_req_1 : boolean;
  signal type_cast_1266_inst_ack_1 : boolean;
  signal type_cast_1276_inst_req_0 : boolean;
  signal type_cast_1276_inst_ack_0 : boolean;
  signal type_cast_1276_inst_req_1 : boolean;
  signal type_cast_1276_inst_ack_1 : boolean;
  signal type_cast_1286_inst_req_0 : boolean;
  signal type_cast_1286_inst_ack_0 : boolean;
  signal type_cast_1286_inst_req_1 : boolean;
  signal type_cast_1286_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1309_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1309_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1309_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1309_inst_ack_1 : boolean;
  signal if_stmt_1323_branch_req_0 : boolean;
  signal if_stmt_1323_branch_ack_1 : boolean;
  signal if_stmt_1323_branch_ack_0 : boolean;
  signal phi_stmt_1195_req_0 : boolean;
  signal type_cast_1201_inst_req_0 : boolean;
  signal type_cast_1201_inst_ack_0 : boolean;
  signal type_cast_1201_inst_req_1 : boolean;
  signal type_cast_1201_inst_ack_1 : boolean;
  signal phi_stmt_1195_req_1 : boolean;
  signal phi_stmt_1195_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_3305_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_3305_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_3305_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_3305_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_3305: Block -- control-path 
    signal sendOutput_CP_3305_elements: BooleanArray(66 downto 0);
    -- 
  begin -- 
    sendOutput_CP_3305_elements(0) <= sendOutput_CP_3305_start;
    sendOutput_CP_3305_symbol <= sendOutput_CP_3305_elements(66);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (83) 
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Sample/word_access_start/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150__entry__
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/branch_block_stmt_1098__entry__
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1098/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/word_access_complete/word_0/$entry
      -- 
    cr_3479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(0), ack => ptr_deref_1133_load_0_req_1); -- 
    cr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(0), ack => ptr_deref_1109_load_0_req_1); -- 
    rr_3468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(0), ack => ptr_deref_1133_load_0_req_0); -- 
    rr_3418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(0), ack => ptr_deref_1121_load_0_req_0); -- 
    rr_3368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(0), ack => ptr_deref_1109_load_0_req_0); -- 
    cr_3429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(0), ack => ptr_deref_1121_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Sample/word_access_start/word_0/ra
      -- 
    ra_3369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_load_0_ack_0, ack => sendOutput_CP_3305_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/ptr_deref_1109_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/ptr_deref_1109_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/ptr_deref_1109_Merge/merge_ack
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/ptr_deref_1109_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1109_Update/word_access_complete/$exit
      -- 
    ca_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_load_0_ack_1, ack => sendOutput_CP_3305_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Sample/word_access_start/word_0/ra
      -- 
    ra_3419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1121_load_0_ack_0, ack => sendOutput_CP_3305_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/ptr_deref_1121_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/ptr_deref_1121_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/ptr_deref_1121_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/ptr_deref_1121_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1121_Update/word_access_complete/word_0/$exit
      -- 
    ca_3430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1121_load_0_ack_1, ack => sendOutput_CP_3305_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Sample/word_access_start/$exit
      -- 
    ra_3469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1133_load_0_ack_0, ack => sendOutput_CP_3305_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/ptr_deref_1133_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/ptr_deref_1133_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/ptr_deref_1133_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_Update/ptr_deref_1133_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/ptr_deref_1133_update_completed_
      -- 
    ca_3480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1133_load_0_ack_1, ack => sendOutput_CP_3305_elements(6)); -- 
    -- CP-element group 7:  branch  join  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (10) 
      -- CP-element group 7: 	 branch_block_stmt_1098/if_stmt_1151_eval_test/$exit
      -- CP-element group 7: 	 branch_block_stmt_1098/if_stmt_1151__entry__
      -- CP-element group 7: 	 branch_block_stmt_1098/R_cmp73_1152_place
      -- CP-element group 7: 	 branch_block_stmt_1098/if_stmt_1151_eval_test/$entry
      -- CP-element group 7: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150/$exit
      -- CP-element group 7: 	 branch_block_stmt_1098/if_stmt_1151_eval_test/branch_req
      -- CP-element group 7: 	 branch_block_stmt_1098/assign_stmt_1106_to_assign_stmt_1150__exit__
      -- CP-element group 7: 	 branch_block_stmt_1098/if_stmt_1151_if_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1098/if_stmt_1151_else_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1098/if_stmt_1151_dead_link/$entry
      -- 
    branch_req_3493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(7), ack => if_stmt_1151_branch_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(2) & sendOutput_CP_3305_elements(4) & sendOutput_CP_3305_elements(6);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (18) 
      -- CP-element group 8: 	 branch_block_stmt_1098/merge_stmt_1157__exit__
      -- CP-element group 8: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192__entry__
      -- CP-element group 8: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/$entry
      -- CP-element group 8: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1098/if_stmt_1151_if_link/$exit
      -- CP-element group 8: 	 branch_block_stmt_1098/if_stmt_1151_if_link/if_choice_transition
      -- CP-element group 8: 	 branch_block_stmt_1098/entry_bbx_xnph
      -- CP-element group 8: 	 branch_block_stmt_1098/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_1098/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 8: 	 branch_block_stmt_1098/merge_stmt_1157_PhiReqMerge
      -- CP-element group 8: 	 branch_block_stmt_1098/merge_stmt_1157_PhiAck/$entry
      -- CP-element group 8: 	 branch_block_stmt_1098/merge_stmt_1157_PhiAck/$exit
      -- CP-element group 8: 	 branch_block_stmt_1098/merge_stmt_1157_PhiAck/dummy
      -- 
    if_choice_transition_3498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1151_branch_ack_1, ack => sendOutput_CP_3305_elements(8)); -- 
    rr_3515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(8), ack => type_cast_1178_inst_req_0); -- 
    cr_3520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(8), ack => type_cast_1178_inst_req_1); -- 
    -- CP-element group 9:  transition  place  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	66 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1098/if_stmt_1151_else_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_1098/entry_forx_xend
      -- CP-element group 9: 	 branch_block_stmt_1098/if_stmt_1151_else_link/else_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_1098/entry_forx_xend_PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_1098/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_3502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1151_branch_ack_0, ack => sendOutput_CP_3305_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_sample_completed_
      -- 
    ra_3516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1178_inst_ack_0, ack => sendOutput_CP_3305_elements(10)); -- 
    -- CP-element group 11:  transition  place  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	60 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192__exit__
      -- CP-element group 11: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody
      -- CP-element group 11: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/$exit
      -- CP-element group 11: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1098/assign_stmt_1163_to_assign_stmt_1192/type_cast_1178_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1195/$entry
      -- CP-element group 11: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/$entry
      -- 
    ca_3521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1178_inst_ack_1, ack => sendOutput_CP_3305_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	65 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	57 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_sample_complete
      -- CP-element group 12: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_Sample/ack
      -- 
    ack_3550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1207_index_offset_ack_0, ack => sendOutput_CP_3305_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	65 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_offset_calculated
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_Update/ack
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_request/req
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_request/$entry
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_Update/$exit
      -- 
    ack_3555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1207_index_offset_ack_1, ack => sendOutput_CP_3305_elements(13)); -- 
    req_3564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(13), ack => addr_of_1208_final_reg_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_request/$exit
      -- CP-element group 14: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_request/ack
      -- 
    ack_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1208_final_reg_ack_0, ack => sendOutput_CP_3305_elements(14)); -- 
    -- CP-element group 15:  join  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	65 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (24) 
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Sample/word_access_start/word_0/rr
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_complete/ack
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_address_resized
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Sample/word_access_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_addr_resize/base_resize_req
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_addr_resize/$entry
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_addr_resize/$exit
      -- CP-element group 15: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_base_addr_resize/base_resize_ack
      -- 
    ack_3570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1208_final_reg_ack_1, ack => sendOutput_CP_3305_elements(15)); -- 
    rr_3603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(15), ack => ptr_deref_1212_load_0_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Sample/word_access_start/word_0/ra
      -- CP-element group 16: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Sample/word_access_start/word_0/$exit
      -- 
    ra_3604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1212_load_0_ack_0, ack => sendOutput_CP_3305_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	65 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	26 
    -- CP-element group 17: 	28 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (33) 
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/ptr_deref_1212_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/ptr_deref_1212_Merge/merge_ack
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/ptr_deref_1212_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/ptr_deref_1212_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_Sample/rr
      -- 
    ca_3615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1212_load_0_ack_1, ack => sendOutput_CP_3305_elements(17)); -- 
    rr_3628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(17), ack => type_cast_1216_inst_req_0); -- 
    rr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(17), ack => type_cast_1226_inst_req_0); -- 
    rr_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(17), ack => type_cast_1236_inst_req_0); -- 
    rr_3670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(17), ack => type_cast_1246_inst_req_0); -- 
    rr_3684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(17), ack => type_cast_1256_inst_req_0); -- 
    rr_3698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(17), ack => type_cast_1266_inst_req_0); -- 
    rr_3712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(17), ack => type_cast_1276_inst_req_0); -- 
    rr_3726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(17), ack => type_cast_1286_inst_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_Sample/$exit
      -- 
    ra_3629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1216_inst_ack_0, ack => sendOutput_CP_3305_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	65 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	54 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_update_completed_
      -- 
    ca_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1216_inst_ack_1, ack => sendOutput_CP_3305_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_Sample/$exit
      -- 
    ra_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1226_inst_ack_0, ack => sendOutput_CP_3305_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	65 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	51 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_update_completed_
      -- 
    ca_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1226_inst_ack_1, ack => sendOutput_CP_3305_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	17 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_Sample/$exit
      -- 
    ra_3657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1236_inst_ack_0, ack => sendOutput_CP_3305_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	65 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	48 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_Update/$exit
      -- 
    ca_3662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1236_inst_ack_1, ack => sendOutput_CP_3305_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_sample_completed_
      -- 
    ra_3671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_0, ack => sendOutput_CP_3305_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	65 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	45 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_update_completed_
      -- 
    ca_3676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_1, ack => sendOutput_CP_3305_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	17 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_Sample/ra
      -- 
    ra_3685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1256_inst_ack_0, ack => sendOutput_CP_3305_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	65 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	42 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_Update/ca
      -- 
    ca_3690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1256_inst_ack_1, ack => sendOutput_CP_3305_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	17 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_Sample/ra
      -- 
    ra_3699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_0, ack => sendOutput_CP_3305_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	65 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	39 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_Update/ca
      -- 
    ca_3704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_1, ack => sendOutput_CP_3305_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_Sample/ra
      -- 
    ra_3713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1276_inst_ack_0, ack => sendOutput_CP_3305_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	65 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_Update/ca
      -- 
    ca_3718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1276_inst_ack_1, ack => sendOutput_CP_3305_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_Sample/ra
      -- 
    ra_3727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1286_inst_ack_0, ack => sendOutput_CP_3305_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	65 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_Sample/req
      -- 
    ca_3732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1286_inst_ack_1, ack => sendOutput_CP_3305_elements(33)); -- 
    req_3740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(33), ack => WPIPE_ConvTranspose_output_pipe_1288_inst_req_0); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_Update/req
      -- 
    ack_3741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0, ack => sendOutput_CP_3305_elements(34)); -- 
    req_3745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(34), ack => WPIPE_ConvTranspose_output_pipe_1288_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1288_Update/ack
      -- 
    ack_3746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1, ack => sendOutput_CP_3305_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	31 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_Sample/req
      -- 
    req_3754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(36), ack => WPIPE_ConvTranspose_output_pipe_1291_inst_req_0); -- 
    sendOutput_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(31) & sendOutput_CP_3305_elements(35);
      gj_sendOutput_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_Update/req
      -- 
    ack_3755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0, ack => sendOutput_CP_3305_elements(37)); -- 
    req_3759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(37), ack => WPIPE_ConvTranspose_output_pipe_1291_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1291_Update/ack
      -- 
    ack_3760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1, ack => sendOutput_CP_3305_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	29 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_Sample/req
      -- 
    req_3768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(39), ack => WPIPE_ConvTranspose_output_pipe_1294_inst_req_0); -- 
    sendOutput_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(29) & sendOutput_CP_3305_elements(38);
      gj_sendOutput_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_Update/req
      -- 
    ack_3769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0, ack => sendOutput_CP_3305_elements(40)); -- 
    req_3773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(40), ack => WPIPE_ConvTranspose_output_pipe_1294_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1294_Update/ack
      -- 
    ack_3774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1, ack => sendOutput_CP_3305_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	27 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_Sample/req
      -- 
    req_3782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(42), ack => WPIPE_ConvTranspose_output_pipe_1297_inst_req_0); -- 
    sendOutput_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(41) & sendOutput_CP_3305_elements(27);
      gj_sendOutput_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_Update/req
      -- 
    ack_3783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0, ack => sendOutput_CP_3305_elements(43)); -- 
    req_3787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(43), ack => WPIPE_ConvTranspose_output_pipe_1297_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1297_Update/ack
      -- 
    ack_3788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1, ack => sendOutput_CP_3305_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	25 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_Sample/req
      -- 
    req_3796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(45), ack => WPIPE_ConvTranspose_output_pipe_1300_inst_req_0); -- 
    sendOutput_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(44) & sendOutput_CP_3305_elements(25);
      gj_sendOutput_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_Update/req
      -- 
    ack_3797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0, ack => sendOutput_CP_3305_elements(46)); -- 
    req_3801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(46), ack => WPIPE_ConvTranspose_output_pipe_1300_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1300_Update/ack
      -- 
    ack_3802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1, ack => sendOutput_CP_3305_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	23 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_Sample/req
      -- 
    req_3810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(48), ack => WPIPE_ConvTranspose_output_pipe_1303_inst_req_0); -- 
    sendOutput_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(47) & sendOutput_CP_3305_elements(23);
      gj_sendOutput_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_Update/req
      -- 
    ack_3811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0, ack => sendOutput_CP_3305_elements(49)); -- 
    req_3815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(49), ack => WPIPE_ConvTranspose_output_pipe_1303_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1303_Update/ack
      -- 
    ack_3816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1, ack => sendOutput_CP_3305_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: 	21 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_Sample/req
      -- 
    req_3824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(51), ack => WPIPE_ConvTranspose_output_pipe_1306_inst_req_0); -- 
    sendOutput_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(50) & sendOutput_CP_3305_elements(21);
      gj_sendOutput_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_Update/req
      -- 
    ack_3825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0, ack => sendOutput_CP_3305_elements(52)); -- 
    req_3829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(52), ack => WPIPE_ConvTranspose_output_pipe_1306_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1306_Update/ack
      -- 
    ack_3830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1, ack => sendOutput_CP_3305_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: 	19 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_Sample/req
      -- 
    req_3838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(54), ack => WPIPE_ConvTranspose_output_pipe_1309_inst_req_0); -- 
    sendOutput_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(53) & sendOutput_CP_3305_elements(19);
      gj_sendOutput_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_Update/req
      -- 
    ack_3839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1309_inst_ack_0, ack => sendOutput_CP_3305_elements(55)); -- 
    req_3843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(55), ack => WPIPE_ConvTranspose_output_pipe_1309_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/WPIPE_ConvTranspose_output_pipe_1309_Update/ack
      -- 
    ack_3844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1309_inst_ack_1, ack => sendOutput_CP_3305_elements(56)); -- 
    -- CP-element group 57:  branch  join  transition  place  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: 	12 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (10) 
      -- CP-element group 57: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322__exit__
      -- CP-element group 57: 	 branch_block_stmt_1098/if_stmt_1323__entry__
      -- CP-element group 57: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/$exit
      -- CP-element group 57: 	 branch_block_stmt_1098/if_stmt_1323_dead_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1098/if_stmt_1323_eval_test/$entry
      -- CP-element group 57: 	 branch_block_stmt_1098/if_stmt_1323_eval_test/$exit
      -- CP-element group 57: 	 branch_block_stmt_1098/if_stmt_1323_eval_test/branch_req
      -- CP-element group 57: 	 branch_block_stmt_1098/R_exitcond1_1324_place
      -- CP-element group 57: 	 branch_block_stmt_1098/if_stmt_1323_if_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1098/if_stmt_1323_else_link/$entry
      -- 
    branch_req_3852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(57), ack => if_stmt_1323_branch_req_0); -- 
    sendOutput_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(56) & sendOutput_CP_3305_elements(12);
      gj_sendOutput_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  merge  transition  place  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	66 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1098/forx_xendx_xloopexit_forx_xend
      -- CP-element group 58: 	 branch_block_stmt_1098/merge_stmt_1329__exit__
      -- CP-element group 58: 	 branch_block_stmt_1098/if_stmt_1323_if_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1098/if_stmt_1323_if_link/if_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1098/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 58: 	 branch_block_stmt_1098/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1098/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1098/merge_stmt_1329_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1098/merge_stmt_1329_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1098/merge_stmt_1329_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1098/merge_stmt_1329_PhiAck/dummy
      -- CP-element group 58: 	 branch_block_stmt_1098/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1098/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1323_branch_ack_1, ack => sendOutput_CP_3305_elements(58)); -- 
    -- CP-element group 59:  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (12) 
      -- CP-element group 59: 	 branch_block_stmt_1098/if_stmt_1323_else_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1098/if_stmt_1323_else_link/else_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/$entry
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/$entry
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1323_branch_ack_0, ack => sendOutput_CP_3305_elements(59)); -- 
    rr_3905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(59), ack => type_cast_1201_inst_req_0); -- 
    cr_3910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(59), ack => type_cast_1201_inst_req_1); -- 
    -- CP-element group 60:  transition  output  delay-element  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	11 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	64 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1195/$exit
      -- CP-element group 60: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/$exit
      -- CP-element group 60: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1199_konst_delay_trans
      -- CP-element group 60: 	 branch_block_stmt_1098/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_req
      -- 
    phi_stmt_1195_req_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1195_req_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(60), ack => phi_stmt_1195_req_0); -- 
    -- Element group sendOutput_CP_3305_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => sendOutput_CP_3305_elements(11), ack => sendOutput_CP_3305_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/Sample/ra
      -- 
    ra_3906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_0, ack => sendOutput_CP_3305_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/Update/ca
      -- 
    ca_3911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_1, ack => sendOutput_CP_3305_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/$exit
      -- CP-element group 63: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/$exit
      -- CP-element group 63: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/$exit
      -- CP-element group 63: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_sources/type_cast_1201/SplitProtocol/$exit
      -- CP-element group 63: 	 branch_block_stmt_1098/forx_xbody_forx_xbody_PhiReq/phi_stmt_1195/phi_stmt_1195_req
      -- 
    phi_stmt_1195_req_3912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1195_req_3912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(63), ack => phi_stmt_1195_req_1); -- 
    sendOutput_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3305_elements(61) & sendOutput_CP_3305_elements(62);
      gj_sendOutput_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3305_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  merge  transition  place  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	60 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1098/merge_stmt_1194_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1098/merge_stmt_1194_PhiAck/$entry
      -- 
    sendOutput_CP_3305_elements(64) <= OrReduce(sendOutput_CP_3305_elements(60) & sendOutput_CP_3305_elements(63));
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	13 
    -- CP-element group 65: 	15 
    -- CP-element group 65: 	17 
    -- CP-element group 65: 	19 
    -- CP-element group 65: 	21 
    -- CP-element group 65: 	23 
    -- CP-element group 65: 	25 
    -- CP-element group 65: 	27 
    -- CP-element group 65: 	29 
    -- CP-element group 65: 	31 
    -- CP-element group 65: 	33 
    -- CP-element group 65:  members (53) 
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_resize_1/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/merge_stmt_1194__exit__
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_resize_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322__entry__
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_scale_1/scale_rename_ack
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_resized_1
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_update_start
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_computed_1
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_scale_1/scale_rename_req
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_Update/req
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/word_access_complete/word_0/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_resize_1/index_resize_ack
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_resize_1/index_resize_req
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1216_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_scale_1/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_complete/req
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/word_access_complete/word_0/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/ptr_deref_1212_Update/word_access_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/addr_of_1208_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_final_index_sum_regn_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1256_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1226_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_scale_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/array_obj_ref_1207_index_scaled_1
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1246_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1236_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1266_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1276_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1098/assign_stmt_1209_to_assign_stmt_1322/type_cast_1286_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1098/merge_stmt_1194_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1098/merge_stmt_1194_PhiAck/phi_stmt_1195_ack
      -- 
    phi_stmt_1195_ack_3917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1195_ack_0, ack => sendOutput_CP_3305_elements(65)); -- 
    req_3554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => array_obj_ref_1207_index_offset_req_1); -- 
    cr_3675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => type_cast_1246_inst_req_1); -- 
    cr_3633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => type_cast_1216_inst_req_1); -- 
    req_3569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => addr_of_1208_final_reg_req_1); -- 
    cr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => type_cast_1226_inst_req_1); -- 
    cr_3614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => ptr_deref_1212_load_0_req_1); -- 
    req_3549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => array_obj_ref_1207_index_offset_req_0); -- 
    cr_3661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => type_cast_1236_inst_req_1); -- 
    cr_3689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => type_cast_1256_inst_req_1); -- 
    cr_3703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => type_cast_1266_inst_req_1); -- 
    cr_3717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => type_cast_1276_inst_req_1); -- 
    cr_3731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3305_elements(65), ack => type_cast_1286_inst_req_1); -- 
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	58 
    -- CP-element group 66: 	9 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 $exit
      -- CP-element group 66: 	 branch_block_stmt_1098/branch_block_stmt_1098__exit__
      -- CP-element group 66: 	 branch_block_stmt_1098/$exit
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1331__exit__
      -- CP-element group 66: 	 branch_block_stmt_1098/return__
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1333__exit__
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1331_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1331_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1331_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1331_PhiAck/dummy
      -- CP-element group 66: 	 branch_block_stmt_1098/return___PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1098/return___PhiReq/$exit
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1333_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1333_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1333_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1098/merge_stmt_1333_PhiAck/dummy
      -- 
    sendOutput_CP_3305_elements(66) <= OrReduce(sendOutput_CP_3305_elements(58) & sendOutput_CP_3305_elements(9));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1206_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1206_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1207_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1209 : std_logic_vector(31 downto 0);
    signal cmp73_1150 : std_logic_vector(0 downto 0);
    signal conv17_1227 : std_logic_vector(7 downto 0);
    signal conv23_1237 : std_logic_vector(7 downto 0);
    signal conv29_1247 : std_logic_vector(7 downto 0);
    signal conv35_1257 : std_logic_vector(7 downto 0);
    signal conv41_1267 : std_logic_vector(7 downto 0);
    signal conv47_1277 : std_logic_vector(7 downto 0);
    signal conv53_1287 : std_logic_vector(7 downto 0);
    signal conv_1217 : std_logic_vector(7 downto 0);
    signal exitcond1_1322 : std_logic_vector(0 downto 0);
    signal iNsTr_0_1106 : std_logic_vector(31 downto 0);
    signal iNsTr_1_1118 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1130 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1179 : std_logic_vector(63 downto 0);
    signal indvar_1195 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1317 : std_logic_vector(63 downto 0);
    signal mul3_1144 : std_logic_vector(31 downto 0);
    signal mul_1139 : std_logic_vector(31 downto 0);
    signal ptr_deref_1109_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1109_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1109_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1109_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1109_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1121_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1121_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1121_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1121_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1121_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1133_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1133_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1133_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1133_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1133_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1212_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1212_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1212_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1212_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1212_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr14_1223 : std_logic_vector(63 downto 0);
    signal shr20_1233 : std_logic_vector(63 downto 0);
    signal shr26_1243 : std_logic_vector(63 downto 0);
    signal shr32_1253 : std_logic_vector(63 downto 0);
    signal shr38_1263 : std_logic_vector(63 downto 0);
    signal shr44_1273 : std_logic_vector(63 downto 0);
    signal shr50_1283 : std_logic_vector(63 downto 0);
    signal tmp1_1122 : std_logic_vector(31 downto 0);
    signal tmp2_1134 : std_logic_vector(31 downto 0);
    signal tmp77_1163 : std_logic_vector(31 downto 0);
    signal tmp77x_xop_1175 : std_logic_vector(31 downto 0);
    signal tmp78_1169 : std_logic_vector(0 downto 0);
    signal tmp81_1192 : std_logic_vector(63 downto 0);
    signal tmp9_1213 : std_logic_vector(63 downto 0);
    signal tmp_1110 : std_logic_vector(31 downto 0);
    signal type_cast_1148_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1161_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1167_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1173_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1183_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1190_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1199_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1201_wire : std_logic_vector(63 downto 0);
    signal type_cast_1221_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1231_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1241_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1251_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1261_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1271_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1281_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1315_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1185 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1207_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1207_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1207_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1207_resized_base_address <= "00000000000000";
    iNsTr_0_1106 <= "00000000000000000000000000000010";
    iNsTr_1_1118 <= "00000000000000000000000000000011";
    iNsTr_2_1130 <= "00000000000000000000000000000100";
    ptr_deref_1109_word_offset_0 <= "0000000";
    ptr_deref_1121_word_offset_0 <= "0000000";
    ptr_deref_1133_word_offset_0 <= "0000000";
    ptr_deref_1212_word_offset_0 <= "00000000000000";
    type_cast_1148_wire_constant <= "00000000000000000000000000000011";
    type_cast_1161_wire_constant <= "00000000000000000000000000000010";
    type_cast_1167_wire_constant <= "00000000000000000000000000000001";
    type_cast_1173_wire_constant <= "11111111111111111111111111111111";
    type_cast_1183_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1190_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1199_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1221_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1231_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1241_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1251_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1261_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1271_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1281_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1315_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1195: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1199_wire_constant & type_cast_1201_wire;
      req <= phi_stmt_1195_req_0 & phi_stmt_1195_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1195",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1195_ack_0,
          idata => idata,
          odata => indvar_1195,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1195
    -- flow-through select operator MUX_1191_inst
    tmp81_1192 <= xx_xop_1185 when (tmp78_1169(0) /=  '0') else type_cast_1190_wire_constant;
    addr_of_1208_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1208_final_reg_req_0;
      addr_of_1208_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1208_final_reg_req_1;
      addr_of_1208_final_reg_ack_1<= rack(0);
      addr_of_1208_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1208_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1207_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1178_inst_req_0;
      type_cast_1178_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1178_inst_req_1;
      type_cast_1178_inst_ack_1<= rack(0);
      type_cast_1178_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1178_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp77x_xop_1175,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_4_1179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1201_inst_req_0;
      type_cast_1201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1201_inst_req_1;
      type_cast_1201_inst_ack_1<= rack(0);
      type_cast_1201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1201_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1216_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1216_inst_req_0;
      type_cast_1216_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1216_inst_req_1;
      type_cast_1216_inst_ack_1<= rack(0);
      type_cast_1216_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1216_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp9_1213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1217,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1226_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1226_inst_req_0;
      type_cast_1226_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1226_inst_req_1;
      type_cast_1226_inst_ack_1<= rack(0);
      type_cast_1226_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1226_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr14_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1227,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1236_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1236_inst_req_0;
      type_cast_1236_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1236_inst_req_1;
      type_cast_1236_inst_ack_1<= rack(0);
      type_cast_1236_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1236_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr20_1233,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_1237,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1246_inst_req_0;
      type_cast_1246_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1246_inst_req_1;
      type_cast_1246_inst_ack_1<= rack(0);
      type_cast_1246_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1246_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr26_1243,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1247,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1256_inst_req_0;
      type_cast_1256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1256_inst_req_1;
      type_cast_1256_inst_ack_1<= rack(0);
      type_cast_1256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr32_1253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_1257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1266_inst_req_0;
      type_cast_1266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1266_inst_req_1;
      type_cast_1266_inst_ack_1<= rack(0);
      type_cast_1266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr38_1263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_1267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1276_inst_req_0;
      type_cast_1276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1276_inst_req_1;
      type_cast_1276_inst_ack_1<= rack(0);
      type_cast_1276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr44_1273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_1277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1286_inst_req_0;
      type_cast_1286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1286_inst_req_1;
      type_cast_1286_inst_ack_1<= rack(0);
      type_cast_1286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr50_1283,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1207_index_1_rename
    process(R_indvar_1206_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1206_resized;
      ov(13 downto 0) := iv;
      R_indvar_1206_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1207_index_1_resize
    process(indvar_1195) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1195;
      ov := iv(13 downto 0);
      R_indvar_1206_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1207_root_address_inst
    process(array_obj_ref_1207_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1207_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1207_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1109_addr_0
    process(ptr_deref_1109_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1109_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1109_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1109_base_resize
    process(iNsTr_0_1106) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_1106;
      ov := iv(6 downto 0);
      ptr_deref_1109_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1109_gather_scatter
    process(ptr_deref_1109_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1109_data_0;
      ov(31 downto 0) := iv;
      tmp_1110 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1109_root_address_inst
    process(ptr_deref_1109_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1109_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1109_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1121_addr_0
    process(ptr_deref_1121_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1121_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1121_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1121_base_resize
    process(iNsTr_1_1118) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_1118;
      ov := iv(6 downto 0);
      ptr_deref_1121_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1121_gather_scatter
    process(ptr_deref_1121_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1121_data_0;
      ov(31 downto 0) := iv;
      tmp1_1122 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1121_root_address_inst
    process(ptr_deref_1121_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1121_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1121_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1133_addr_0
    process(ptr_deref_1133_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1133_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1133_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1133_base_resize
    process(iNsTr_2_1130) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1130;
      ov := iv(6 downto 0);
      ptr_deref_1133_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1133_gather_scatter
    process(ptr_deref_1133_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1133_data_0;
      ov(31 downto 0) := iv;
      tmp2_1134 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1133_root_address_inst
    process(ptr_deref_1133_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1133_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1133_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1212_addr_0
    process(ptr_deref_1212_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1212_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1212_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1212_base_resize
    process(arrayidx_1209) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1209;
      ov := iv(13 downto 0);
      ptr_deref_1212_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1212_gather_scatter
    process(ptr_deref_1212_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1212_data_0;
      ov(63 downto 0) := iv;
      tmp9_1213 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1212_root_address_inst
    process(ptr_deref_1212_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1212_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1212_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1151_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp73_1150;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1151_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1151_branch_req_0,
          ack0 => if_stmt_1151_branch_ack_0,
          ack1 => if_stmt_1151_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1323_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1322;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1323_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1323_branch_req_0,
          ack0 => if_stmt_1323_branch_ack_0,
          ack1 => if_stmt_1323_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1174_inst
    process(tmp77_1163) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp77_1163, type_cast_1173_wire_constant, tmp_var);
      tmp77x_xop_1175 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1184_inst
    process(iNsTr_4_1179) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_4_1179, type_cast_1183_wire_constant, tmp_var);
      xx_xop_1185 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1316_inst
    process(indvar_1195) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1195, type_cast_1315_wire_constant, tmp_var);
      indvarx_xnext_1317 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1321_inst
    process(indvarx_xnext_1317, tmp81_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1317, tmp81_1192, tmp_var);
      exitcond1_1322 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1162_inst
    process(mul3_1144) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul3_1144, type_cast_1161_wire_constant, tmp_var);
      tmp77_1163 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1222_inst
    process(tmp9_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1213, type_cast_1221_wire_constant, tmp_var);
      shr14_1223 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1232_inst
    process(tmp9_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1213, type_cast_1231_wire_constant, tmp_var);
      shr20_1233 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1242_inst
    process(tmp9_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1213, type_cast_1241_wire_constant, tmp_var);
      shr26_1243 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1252_inst
    process(tmp9_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1213, type_cast_1251_wire_constant, tmp_var);
      shr32_1253 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1262_inst
    process(tmp9_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1213, type_cast_1261_wire_constant, tmp_var);
      shr38_1263 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1272_inst
    process(tmp9_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1213, type_cast_1271_wire_constant, tmp_var);
      shr44_1273 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1282_inst
    process(tmp9_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1213, type_cast_1281_wire_constant, tmp_var);
      shr50_1283 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1138_inst
    process(tmp1_1122, tmp_1110) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1122, tmp_1110, tmp_var);
      mul_1139 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1143_inst
    process(mul_1139, tmp2_1134) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1139, tmp2_1134, tmp_var);
      mul3_1144 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1149_inst
    process(mul3_1144) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul3_1144, type_cast_1148_wire_constant, tmp_var);
      cmp73_1150 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1168_inst
    process(tmp77_1163) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp77_1163, type_cast_1167_wire_constant, tmp_var);
      tmp78_1169 <= tmp_var; --
    end process;
    -- shared split operator group (16) : array_obj_ref_1207_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1206_scaled;
      array_obj_ref_1207_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1207_index_offset_req_0;
      array_obj_ref_1207_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1207_index_offset_req_1;
      array_obj_ref_1207_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared load operator group (0) : ptr_deref_1133_load_0 ptr_deref_1121_load_0 ptr_deref_1109_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1133_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1121_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1109_load_0_req_0;
      ptr_deref_1133_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1121_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1109_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1133_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1121_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1109_load_0_req_1;
      ptr_deref_1133_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1121_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1109_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1133_word_address_0 & ptr_deref_1121_word_address_0 & ptr_deref_1109_word_address_0;
      ptr_deref_1133_data_0 <= data_out(95 downto 64);
      ptr_deref_1121_data_0 <= data_out(63 downto 32);
      ptr_deref_1109_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1212_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1212_load_0_req_0;
      ptr_deref_1212_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1212_load_0_req_1;
      ptr_deref_1212_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1212_word_address_0;
      ptr_deref_1212_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(13 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(63 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1291_inst WPIPE_ConvTranspose_output_pipe_1288_inst WPIPE_ConvTranspose_output_pipe_1306_inst WPIPE_ConvTranspose_output_pipe_1309_inst WPIPE_ConvTranspose_output_pipe_1303_inst WPIPE_ConvTranspose_output_pipe_1300_inst WPIPE_ConvTranspose_output_pipe_1297_inst WPIPE_ConvTranspose_output_pipe_1294_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1291_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1288_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1306_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1309_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1303_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1300_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1297_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1294_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1309_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1291_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1288_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1306_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1309_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1303_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1300_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1297_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1294_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1309_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv47_1277 & conv53_1287 & conv17_1227 & conv_1217 & conv23_1237 & conv29_1247 & conv35_1257 & conv41_1267;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_0_start: Boolean;
  signal testConfigure_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_469_load_0_ack_0 : boolean;
  signal ptr_deref_383_load_0_req_0 : boolean;
  signal type_cast_898_inst_req_1 : boolean;
  signal ptr_deref_469_load_0_req_0 : boolean;
  signal ptr_deref_469_load_0_ack_1 : boolean;
  signal type_cast_916_inst_ack_1 : boolean;
  signal if_stmt_502_branch_ack_1 : boolean;
  signal if_stmt_502_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_ack_0 : boolean;
  signal if_stmt_502_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_36_inst_ack_1 : boolean;
  signal ptr_deref_370_store_0_ack_1 : boolean;
  signal ptr_deref_370_store_0_req_1 : boolean;
  signal type_cast_359_inst_ack_0 : boolean;
  signal ptr_deref_370_store_0_ack_0 : boolean;
  signal ptr_deref_370_store_0_req_0 : boolean;
  signal type_cast_880_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_36_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_36_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_36_inst_req_1 : boolean;
  signal ptr_deref_433_load_0_ack_0 : boolean;
  signal ptr_deref_433_load_0_req_0 : boolean;
  signal type_cast_359_inst_ack_1 : boolean;
  signal type_cast_40_inst_req_0 : boolean;
  signal type_cast_40_inst_ack_0 : boolean;
  signal type_cast_40_inst_req_1 : boolean;
  signal type_cast_40_inst_ack_1 : boolean;
  signal type_cast_488_inst_req_1 : boolean;
  signal ptr_deref_457_load_0_ack_1 : boolean;
  signal ptr_deref_957_load_0_ack_0 : boolean;
  signal ptr_deref_457_load_0_req_1 : boolean;
  signal ptr_deref_49_store_0_req_0 : boolean;
  signal ptr_deref_49_store_0_ack_0 : boolean;
  signal ptr_deref_49_store_0_req_1 : boolean;
  signal ptr_deref_49_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal ptr_deref_445_load_0_ack_1 : boolean;
  signal if_stmt_66_branch_req_0 : boolean;
  signal if_stmt_66_branch_ack_1 : boolean;
  signal ptr_deref_407_load_0_ack_1 : boolean;
  signal if_stmt_66_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_req_0 : boolean;
  signal ptr_deref_407_load_0_req_1 : boolean;
  signal ptr_deref_445_load_0_req_1 : boolean;
  signal type_cast_97_inst_req_0 : boolean;
  signal type_cast_97_inst_ack_0 : boolean;
  signal type_cast_97_inst_req_1 : boolean;
  signal type_cast_97_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_ack_1 : boolean;
  signal type_cast_488_inst_ack_0 : boolean;
  signal ptr_deref_433_load_0_ack_1 : boolean;
  signal ptr_deref_433_load_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_ack_0 : boolean;
  signal array_obj_ref_103_index_offset_req_0 : boolean;
  signal array_obj_ref_103_index_offset_ack_0 : boolean;
  signal array_obj_ref_103_index_offset_req_1 : boolean;
  signal array_obj_ref_103_index_offset_ack_1 : boolean;
  signal ptr_deref_981_load_0_req_0 : boolean;
  signal addr_of_104_final_reg_req_0 : boolean;
  signal addr_of_104_final_reg_ack_0 : boolean;
  signal addr_of_104_final_reg_req_1 : boolean;
  signal addr_of_104_final_reg_ack_1 : boolean;
  signal type_cast_488_inst_req_0 : boolean;
  signal ptr_deref_981_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_ack_0 : boolean;
  signal ptr_deref_981_load_0_req_1 : boolean;
  signal ptr_deref_107_store_0_req_0 : boolean;
  signal ptr_deref_107_store_0_ack_0 : boolean;
  signal ptr_deref_457_load_0_ack_0 : boolean;
  signal ptr_deref_107_store_0_req_1 : boolean;
  signal ptr_deref_107_store_0_ack_1 : boolean;
  signal ptr_deref_395_load_0_ack_1 : boolean;
  signal addr_of_276_final_reg_req_0 : boolean;
  signal addr_of_276_final_reg_ack_0 : boolean;
  signal addr_of_276_final_reg_req_1 : boolean;
  signal addr_of_276_final_reg_ack_1 : boolean;
  signal ptr_deref_395_load_0_req_1 : boolean;
  signal ptr_deref_457_load_0_req_0 : boolean;
  signal type_cast_421_inst_ack_1 : boolean;
  signal ptr_deref_124_load_0_req_0 : boolean;
  signal ptr_deref_124_load_0_ack_0 : boolean;
  signal ptr_deref_124_load_0_req_1 : boolean;
  signal ptr_deref_124_load_0_ack_1 : boolean;
  signal if_stmt_999_branch_req_0 : boolean;
  signal type_cast_359_inst_req_1 : boolean;
  signal type_cast_1026_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_132_inst_req_0 : boolean;
  signal type_cast_421_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_132_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_132_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_132_inst_ack_1 : boolean;
  signal type_cast_136_inst_req_0 : boolean;
  signal type_cast_136_inst_ack_0 : boolean;
  signal type_cast_136_inst_req_1 : boolean;
  signal type_cast_136_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_req_1 : boolean;
  signal ptr_deref_445_load_0_ack_0 : boolean;
  signal if_stmt_138_branch_req_0 : boolean;
  signal if_stmt_138_branch_ack_1 : boolean;
  signal if_stmt_138_branch_ack_0 : boolean;
  signal type_cast_1026_inst_ack_0 : boolean;
  signal type_cast_421_inst_ack_0 : boolean;
  signal ptr_deref_445_load_0_req_0 : boolean;
  signal type_cast_421_inst_req_0 : boolean;
  signal ptr_deref_166_store_0_req_0 : boolean;
  signal ptr_deref_166_store_0_ack_0 : boolean;
  signal ptr_deref_166_store_0_req_1 : boolean;
  signal ptr_deref_166_store_0_ack_1 : boolean;
  signal ptr_deref_407_load_0_ack_0 : boolean;
  signal if_stmt_175_branch_req_0 : boolean;
  signal if_stmt_175_branch_ack_1 : boolean;
  signal ptr_deref_407_load_0_req_0 : boolean;
  signal if_stmt_175_branch_ack_0 : boolean;
  signal type_cast_200_inst_req_0 : boolean;
  signal type_cast_200_inst_ack_0 : boolean;
  signal type_cast_200_inst_req_1 : boolean;
  signal type_cast_200_inst_ack_1 : boolean;
  signal array_obj_ref_206_index_offset_req_0 : boolean;
  signal array_obj_ref_206_index_offset_ack_0 : boolean;
  signal array_obj_ref_206_index_offset_req_1 : boolean;
  signal array_obj_ref_206_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_ack_1 : boolean;
  signal addr_of_207_final_reg_req_0 : boolean;
  signal addr_of_207_final_reg_ack_0 : boolean;
  signal addr_of_207_final_reg_req_1 : boolean;
  signal ptr_deref_957_load_0_req_0 : boolean;
  signal addr_of_207_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_210_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_210_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_210_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_210_inst_ack_1 : boolean;
  signal type_cast_214_inst_req_0 : boolean;
  signal type_cast_214_inst_ack_0 : boolean;
  signal type_cast_214_inst_req_1 : boolean;
  signal type_cast_214_inst_ack_1 : boolean;
  signal ptr_deref_383_load_0_ack_1 : boolean;
  signal ptr_deref_383_load_0_req_1 : boolean;
  signal ptr_deref_217_store_0_req_0 : boolean;
  signal ptr_deref_217_store_0_ack_0 : boolean;
  signal ptr_deref_217_store_0_req_1 : boolean;
  signal ptr_deref_217_store_0_ack_1 : boolean;
  signal if_stmt_999_branch_ack_1 : boolean;
  signal ptr_deref_234_load_0_req_0 : boolean;
  signal ptr_deref_234_load_0_ack_0 : boolean;
  signal ptr_deref_234_load_0_req_1 : boolean;
  signal ptr_deref_234_load_0_ack_1 : boolean;
  signal type_cast_488_inst_ack_1 : boolean;
  signal type_cast_898_inst_ack_1 : boolean;
  signal ptr_deref_469_load_0_req_1 : boolean;
  signal if_stmt_241_branch_req_0 : boolean;
  signal if_stmt_241_branch_ack_1 : boolean;
  signal type_cast_359_inst_req_0 : boolean;
  signal if_stmt_241_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_251_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_251_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_251_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_251_inst_ack_1 : boolean;
  signal ptr_deref_957_load_0_req_1 : boolean;
  signal type_cast_255_inst_req_0 : boolean;
  signal type_cast_255_inst_ack_0 : boolean;
  signal type_cast_255_inst_req_1 : boolean;
  signal type_cast_255_inst_ack_1 : boolean;
  signal ptr_deref_395_load_0_ack_0 : boolean;
  signal ptr_deref_395_load_0_req_0 : boolean;
  signal ptr_deref_383_load_0_ack_0 : boolean;
  signal ptr_deref_279_store_0_req_0 : boolean;
  signal ptr_deref_279_store_0_ack_0 : boolean;
  signal ptr_deref_957_load_0_ack_1 : boolean;
  signal ptr_deref_279_store_0_req_1 : boolean;
  signal ptr_deref_279_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_283_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_283_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_283_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_283_inst_ack_1 : boolean;
  signal type_cast_862_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_req_1 : boolean;
  signal type_cast_287_inst_req_0 : boolean;
  signal type_cast_287_inst_ack_0 : boolean;
  signal type_cast_287_inst_req_1 : boolean;
  signal type_cast_287_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_ack_1 : boolean;
  signal type_cast_862_inst_ack_0 : boolean;
  signal if_stmt_301_branch_req_0 : boolean;
  signal ptr_deref_969_load_0_req_0 : boolean;
  signal if_stmt_301_branch_ack_1 : boolean;
  signal if_stmt_301_branch_ack_0 : boolean;
  signal ptr_deref_969_load_0_ack_0 : boolean;
  signal type_cast_880_inst_req_0 : boolean;
  signal STORE_padding_313_store_0_req_0 : boolean;
  signal STORE_padding_313_store_0_ack_0 : boolean;
  signal STORE_padding_313_store_0_req_1 : boolean;
  signal STORE_padding_313_store_0_ack_1 : boolean;
  signal if_stmt_999_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_317_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_317_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_317_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_317_inst_ack_1 : boolean;
  signal type_cast_862_inst_req_1 : boolean;
  signal type_cast_862_inst_ack_1 : boolean;
  signal type_cast_321_inst_req_0 : boolean;
  signal type_cast_321_inst_ack_0 : boolean;
  signal type_cast_321_inst_req_1 : boolean;
  signal type_cast_321_inst_ack_1 : boolean;
  signal ptr_deref_332_store_0_req_0 : boolean;
  signal ptr_deref_332_store_0_ack_0 : boolean;
  signal ptr_deref_332_store_0_req_1 : boolean;
  signal ptr_deref_332_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_ack_1 : boolean;
  signal type_cast_340_inst_req_0 : boolean;
  signal type_cast_340_inst_ack_0 : boolean;
  signal type_cast_340_inst_req_1 : boolean;
  signal type_cast_340_inst_ack_1 : boolean;
  signal ptr_deref_351_store_0_req_0 : boolean;
  signal ptr_deref_351_store_0_ack_0 : boolean;
  signal ptr_deref_351_store_0_req_1 : boolean;
  signal ptr_deref_351_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_355_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_355_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_355_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_355_inst_ack_1 : boolean;
  signal type_cast_916_inst_req_1 : boolean;
  signal if_stmt_523_branch_req_0 : boolean;
  signal if_stmt_523_branch_ack_1 : boolean;
  signal if_stmt_523_branch_ack_0 : boolean;
  signal type_cast_542_inst_req_0 : boolean;
  signal type_cast_542_inst_ack_0 : boolean;
  signal type_cast_542_inst_req_1 : boolean;
  signal type_cast_542_inst_ack_1 : boolean;
  signal ptr_deref_1059_store_0_req_0 : boolean;
  signal type_cast_1026_inst_ack_1 : boolean;
  signal array_obj_ref_577_index_offset_req_0 : boolean;
  signal array_obj_ref_577_index_offset_ack_0 : boolean;
  signal type_cast_898_inst_ack_0 : boolean;
  signal array_obj_ref_577_index_offset_req_1 : boolean;
  signal array_obj_ref_577_index_offset_ack_1 : boolean;
  signal type_cast_898_inst_req_0 : boolean;
  signal addr_of_578_final_reg_req_0 : boolean;
  signal addr_of_578_final_reg_ack_0 : boolean;
  signal addr_of_578_final_reg_req_1 : boolean;
  signal addr_of_578_final_reg_ack_1 : boolean;
  signal addr_of_1056_final_reg_ack_1 : boolean;
  signal if_stmt_938_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_581_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_581_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_581_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_581_inst_ack_1 : boolean;
  signal array_obj_ref_1055_index_offset_ack_1 : boolean;
  signal type_cast_585_inst_req_0 : boolean;
  signal type_cast_585_inst_ack_0 : boolean;
  signal type_cast_585_inst_req_1 : boolean;
  signal type_cast_585_inst_ack_1 : boolean;
  signal addr_of_1056_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_594_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_594_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_594_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_594_inst_ack_1 : boolean;
  signal array_obj_ref_1055_index_offset_req_1 : boolean;
  signal if_stmt_938_branch_ack_1 : boolean;
  signal type_cast_598_inst_req_0 : boolean;
  signal type_cast_598_inst_ack_0 : boolean;
  signal type_cast_598_inst_req_1 : boolean;
  signal type_cast_598_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_612_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_612_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_612_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_612_inst_ack_1 : boolean;
  signal if_stmt_938_branch_req_0 : boolean;
  signal type_cast_616_inst_req_0 : boolean;
  signal type_cast_616_inst_ack_0 : boolean;
  signal type_cast_616_inst_req_1 : boolean;
  signal type_cast_616_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_630_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_630_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_630_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_630_inst_ack_1 : boolean;
  signal type_cast_634_inst_req_0 : boolean;
  signal type_cast_634_inst_ack_0 : boolean;
  signal type_cast_634_inst_req_1 : boolean;
  signal type_cast_634_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_648_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_648_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_648_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_648_inst_ack_1 : boolean;
  signal array_obj_ref_1055_index_offset_ack_0 : boolean;
  signal array_obj_ref_1055_index_offset_req_0 : boolean;
  signal type_cast_652_inst_req_0 : boolean;
  signal type_cast_652_inst_ack_0 : boolean;
  signal type_cast_652_inst_req_1 : boolean;
  signal type_cast_652_inst_ack_1 : boolean;
  signal addr_of_1056_final_reg_ack_0 : boolean;
  signal type_cast_844_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_666_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_666_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_666_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_666_inst_ack_1 : boolean;
  signal ptr_deref_924_store_0_ack_1 : boolean;
  signal type_cast_670_inst_req_0 : boolean;
  signal type_cast_670_inst_ack_0 : boolean;
  signal type_cast_670_inst_req_1 : boolean;
  signal type_cast_670_inst_ack_1 : boolean;
  signal addr_of_1056_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_684_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_684_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_684_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_684_inst_ack_1 : boolean;
  signal ptr_deref_924_store_0_req_1 : boolean;
  signal type_cast_688_inst_req_0 : boolean;
  signal type_cast_688_inst_ack_0 : boolean;
  signal type_cast_688_inst_req_1 : boolean;
  signal type_cast_688_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_702_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_702_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_702_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_702_inst_ack_1 : boolean;
  signal type_cast_1026_inst_req_1 : boolean;
  signal type_cast_706_inst_req_0 : boolean;
  signal ptr_deref_969_load_0_ack_1 : boolean;
  signal type_cast_706_inst_ack_0 : boolean;
  signal type_cast_706_inst_req_1 : boolean;
  signal ptr_deref_969_load_0_req_1 : boolean;
  signal type_cast_706_inst_ack_1 : boolean;
  signal ptr_deref_1059_store_0_ack_0 : boolean;
  signal ptr_deref_981_load_0_ack_1 : boolean;
  signal ptr_deref_924_store_0_ack_0 : boolean;
  signal ptr_deref_924_store_0_req_0 : boolean;
  signal type_cast_916_inst_ack_0 : boolean;
  signal ptr_deref_714_store_0_req_0 : boolean;
  signal ptr_deref_714_store_0_ack_0 : boolean;
  signal type_cast_844_inst_req_1 : boolean;
  signal type_cast_916_inst_req_0 : boolean;
  signal ptr_deref_714_store_0_req_1 : boolean;
  signal ptr_deref_714_store_0_ack_1 : boolean;
  signal type_cast_880_inst_ack_1 : boolean;
  signal type_cast_880_inst_req_1 : boolean;
  signal if_stmt_728_branch_req_0 : boolean;
  signal if_stmt_728_branch_ack_1 : boolean;
  signal if_stmt_728_branch_ack_0 : boolean;
  signal type_cast_752_inst_req_0 : boolean;
  signal type_cast_752_inst_ack_0 : boolean;
  signal type_cast_752_inst_req_1 : boolean;
  signal type_cast_752_inst_ack_1 : boolean;
  signal array_obj_ref_787_index_offset_req_0 : boolean;
  signal array_obj_ref_787_index_offset_ack_0 : boolean;
  signal array_obj_ref_787_index_offset_req_1 : boolean;
  signal array_obj_ref_787_index_offset_ack_1 : boolean;
  signal addr_of_788_final_reg_req_0 : boolean;
  signal addr_of_788_final_reg_ack_0 : boolean;
  signal addr_of_788_final_reg_req_1 : boolean;
  signal addr_of_788_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_791_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_791_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_791_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_791_inst_ack_1 : boolean;
  signal type_cast_795_inst_req_0 : boolean;
  signal type_cast_795_inst_ack_0 : boolean;
  signal type_cast_795_inst_req_1 : boolean;
  signal type_cast_795_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_804_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_804_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_804_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_804_inst_ack_1 : boolean;
  signal type_cast_808_inst_req_0 : boolean;
  signal type_cast_808_inst_ack_0 : boolean;
  signal type_cast_808_inst_req_1 : boolean;
  signal type_cast_808_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_822_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_822_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_822_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_822_inst_ack_1 : boolean;
  signal type_cast_826_inst_req_0 : boolean;
  signal type_cast_826_inst_ack_0 : boolean;
  signal type_cast_826_inst_req_1 : boolean;
  signal type_cast_826_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_840_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_840_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_840_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_840_inst_ack_1 : boolean;
  signal type_cast_844_inst_req_0 : boolean;
  signal type_cast_844_inst_ack_0 : boolean;
  signal ptr_deref_1059_store_0_req_1 : boolean;
  signal ptr_deref_1059_store_0_ack_1 : boolean;
  signal if_stmt_1074_branch_req_0 : boolean;
  signal if_stmt_1074_branch_ack_1 : boolean;
  signal if_stmt_1074_branch_ack_0 : boolean;
  signal type_cast_1085_inst_req_0 : boolean;
  signal type_cast_1085_inst_ack_0 : boolean;
  signal type_cast_1085_inst_req_1 : boolean;
  signal type_cast_1085_inst_ack_1 : boolean;
  signal type_cast_78_inst_req_0 : boolean;
  signal type_cast_78_inst_ack_0 : boolean;
  signal type_cast_78_inst_req_1 : boolean;
  signal type_cast_78_inst_ack_1 : boolean;
  signal phi_stmt_75_req_0 : boolean;
  signal type_cast_85_inst_req_0 : boolean;
  signal type_cast_85_inst_ack_0 : boolean;
  signal type_cast_85_inst_req_1 : boolean;
  signal type_cast_85_inst_ack_1 : boolean;
  signal phi_stmt_82_req_0 : boolean;
  signal phi_stmt_75_req_1 : boolean;
  signal type_cast_87_inst_req_0 : boolean;
  signal type_cast_87_inst_ack_0 : boolean;
  signal type_cast_87_inst_req_1 : boolean;
  signal type_cast_87_inst_ack_1 : boolean;
  signal phi_stmt_82_req_1 : boolean;
  signal phi_stmt_75_ack_0 : boolean;
  signal phi_stmt_82_ack_0 : boolean;
  signal type_cast_148_inst_req_0 : boolean;
  signal type_cast_148_inst_ack_0 : boolean;
  signal type_cast_148_inst_req_1 : boolean;
  signal type_cast_148_inst_ack_1 : boolean;
  signal phi_stmt_145_req_0 : boolean;
  signal phi_stmt_145_ack_0 : boolean;
  signal type_cast_155_inst_req_0 : boolean;
  signal type_cast_155_inst_ack_0 : boolean;
  signal type_cast_155_inst_req_1 : boolean;
  signal type_cast_155_inst_ack_1 : boolean;
  signal phi_stmt_152_req_0 : boolean;
  signal type_cast_157_inst_req_0 : boolean;
  signal type_cast_157_inst_ack_0 : boolean;
  signal type_cast_157_inst_req_1 : boolean;
  signal type_cast_157_inst_ack_1 : boolean;
  signal phi_stmt_152_req_1 : boolean;
  signal phi_stmt_152_ack_0 : boolean;
  signal type_cast_187_inst_req_0 : boolean;
  signal type_cast_187_inst_ack_0 : boolean;
  signal type_cast_187_inst_req_1 : boolean;
  signal type_cast_187_inst_ack_1 : boolean;
  signal phi_stmt_184_req_0 : boolean;
  signal phi_stmt_184_req_1 : boolean;
  signal phi_stmt_184_ack_0 : boolean;
  signal phi_stmt_259_req_0 : boolean;
  signal type_cast_269_inst_req_0 : boolean;
  signal type_cast_269_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_1 : boolean;
  signal type_cast_269_inst_ack_1 : boolean;
  signal phi_stmt_266_req_0 : boolean;
  signal type_cast_265_inst_req_0 : boolean;
  signal type_cast_265_inst_ack_0 : boolean;
  signal type_cast_265_inst_req_1 : boolean;
  signal type_cast_265_inst_ack_1 : boolean;
  signal phi_stmt_259_req_1 : boolean;
  signal type_cast_271_inst_req_0 : boolean;
  signal type_cast_271_inst_ack_0 : boolean;
  signal type_cast_271_inst_req_1 : boolean;
  signal type_cast_271_inst_ack_1 : boolean;
  signal phi_stmt_266_req_1 : boolean;
  signal phi_stmt_259_ack_0 : boolean;
  signal phi_stmt_266_ack_0 : boolean;
  signal type_cast_311_inst_req_0 : boolean;
  signal type_cast_311_inst_ack_0 : boolean;
  signal type_cast_311_inst_req_1 : boolean;
  signal type_cast_311_inst_ack_1 : boolean;
  signal phi_stmt_308_req_0 : boolean;
  signal phi_stmt_308_ack_0 : boolean;
  signal phi_stmt_565_req_0 : boolean;
  signal type_cast_571_inst_req_0 : boolean;
  signal type_cast_571_inst_ack_0 : boolean;
  signal type_cast_571_inst_req_1 : boolean;
  signal type_cast_571_inst_ack_1 : boolean;
  signal phi_stmt_565_req_1 : boolean;
  signal phi_stmt_565_ack_0 : boolean;
  signal phi_stmt_775_req_0 : boolean;
  signal type_cast_781_inst_req_0 : boolean;
  signal type_cast_781_inst_ack_0 : boolean;
  signal type_cast_781_inst_req_1 : boolean;
  signal type_cast_781_inst_ack_1 : boolean;
  signal phi_stmt_775_req_1 : boolean;
  signal phi_stmt_775_ack_0 : boolean;
  signal phi_stmt_1043_req_0 : boolean;
  signal type_cast_1049_inst_req_0 : boolean;
  signal type_cast_1049_inst_ack_0 : boolean;
  signal type_cast_1049_inst_req_1 : boolean;
  signal type_cast_1049_inst_ack_1 : boolean;
  signal phi_stmt_1043_req_1 : boolean;
  signal phi_stmt_1043_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_0: Block -- control-path 
    signal testConfigure_CP_0_elements: BooleanArray(310 downto 0);
    -- 
  begin -- 
    testConfigure_CP_0_elements(0) <= testConfigure_CP_0_start;
    testConfigure_CP_0_symbol <= testConfigure_CP_0_elements(233);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (35) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_34/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/branch_block_stmt_34__entry__
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65__entry__
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_update_start_
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_Update/cr
      -- 
    rr_118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => RPIPE_ConvTranspose_input_pipe_36_inst_req_0); -- 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_40_inst_req_1); -- 
    cr_187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => ptr_deref_49_store_0_req_1); -- 
    cr_215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_64_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_update_start_
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_Update/cr
      -- 
    ra_119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_36_inst_ack_0, ack => testConfigure_CP_0_elements(1)); -- 
    cr_123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(1), ack => RPIPE_ConvTranspose_input_pipe_36_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_36_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_Sample/rr
      -- 
    ca_124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_36_inst_ack_1, ack => testConfigure_CP_0_elements(2)); -- 
    rr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => type_cast_40_inst_req_0); -- 
    rr_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_Sample/ra
      -- 
    ra_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_40_inst_ack_0, ack => testConfigure_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_40_Update/ca
      -- 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_40_inst_ack_1, ack => testConfigure_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/ptr_deref_49_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/ptr_deref_49_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/ptr_deref_49_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/ptr_deref_49_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/word_access_start/word_0/rr
      -- 
    rr_176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(5), ack => ptr_deref_49_store_0_req_0); -- 
    testConfigure_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(0) & testConfigure_CP_0_elements(4);
      gj_testConfigure_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Sample/word_access_start/word_0/ra
      -- 
    ra_177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_49_store_0_ack_0, ack => testConfigure_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/ptr_deref_49_Update/word_access_complete/word_0/ca
      -- 
    ca_188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_49_store_0_ack_1, ack => testConfigure_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_update_start_
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_Update/cr
      -- 
    ra_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_0, ack => testConfigure_CP_0_elements(8)); -- 
    cr_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(8), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/RPIPE_ConvTranspose_input_pipe_60_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_Sample/rr
      -- 
    ca_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_1, ack => testConfigure_CP_0_elements(9)); -- 
    rr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(9), ack => type_cast_64_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_Sample/ra
      -- 
    ra_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => testConfigure_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/type_cast_64_Update/ca
      -- 
    ca_216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => testConfigure_CP_0_elements(11)); -- 
    -- CP-element group 12:  branch  join  transition  place  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (10) 
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65__exit__
      -- CP-element group 12: 	 branch_block_stmt_34/if_stmt_66__entry__
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_37_to_assign_stmt_65/$exit
      -- CP-element group 12: 	 branch_block_stmt_34/if_stmt_66_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_34/if_stmt_66_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_34/if_stmt_66_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_34/if_stmt_66_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_34/R_cmp227_67_place
      -- CP-element group 12: 	 branch_block_stmt_34/if_stmt_66_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_34/if_stmt_66_else_link/$entry
      -- 
    branch_req_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(12), ack => if_stmt_66_branch_req_0); -- 
    testConfigure_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(7) & testConfigure_CP_0_elements(11);
      gj_testConfigure_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	254 
    -- CP-element group 13: 	255 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_34/if_stmt_66_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_34/if_stmt_66_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/Update/cr
      -- 
    if_choice_transition_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_66_branch_ack_1, ack => testConfigure_CP_0_elements(13)); -- 
    rr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_155_inst_req_0); -- 
    cr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_155_inst_req_1); -- 
    -- CP-element group 14:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	241 
    -- CP-element group 14: 	242 
    -- CP-element group 14: 	243 
    -- CP-element group 14:  members (22) 
      -- CP-element group 14: 	 branch_block_stmt_34/merge_stmt_72__exit__
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 14: 	 branch_block_stmt_34/if_stmt_66_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_34/if_stmt_66_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_34/entry_forx_xbodyx_xpreheader
      -- CP-element group 14: 	 branch_block_stmt_34/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_34/merge_stmt_72_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_34/merge_stmt_72_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/merge_stmt_72_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_34/merge_stmt_72_PhiAck/dummy
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_75/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/Update/cr
      -- 
    else_choice_transition_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_66_branch_ack_0, ack => testConfigure_CP_0_elements(14)); -- 
    rr_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_87_inst_req_0); -- 
    cr_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_87_inst_req_1); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	249 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_Sample/ra
      -- 
    ra_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_97_inst_ack_0, ack => testConfigure_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	249 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_Update/ca
      -- 
    ca_252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_97_inst_ack_1, ack => testConfigure_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	249 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	31 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_sample_complete
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_Sample/ack
      -- 
    ack_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_103_index_offset_ack_0, ack => testConfigure_CP_0_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	249 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (11) 
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_Update/ack
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_request/$entry
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_request/req
      -- 
    ack_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_103_index_offset_ack_1, ack => testConfigure_CP_0_elements(18)); -- 
    req_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(18), ack => addr_of_104_final_reg_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_request/$exit
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_request/ack
      -- 
    ack_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_104_final_reg_ack_0, ack => testConfigure_CP_0_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	249 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (28) 
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_complete/ack
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_word_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_root_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_address_resized
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_addr_resize/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_addr_resize/$exit
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_addr_resize/base_resize_req
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_addr_resize/base_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_plus_offset/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_plus_offset/$exit
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_plus_offset/sum_rename_req
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_base_plus_offset/sum_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_word_addrgen/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_word_addrgen/$exit
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_word_addrgen/root_register_req
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_word_addrgen/root_register_ack
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/ptr_deref_107_Split/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/ptr_deref_107_Split/$exit
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/ptr_deref_107_Split/split_req
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/ptr_deref_107_Split/split_ack
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/word_access_start/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/word_access_start/word_0/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/word_access_start/word_0/rr
      -- 
    ack_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_104_final_reg_ack_1, ack => testConfigure_CP_0_elements(20)); -- 
    rr_336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(20), ack => ptr_deref_107_store_0_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	30 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Sample/word_access_start/word_0/ra
      -- 
    ra_337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_107_store_0_ack_0, ack => testConfigure_CP_0_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	249 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Update/word_access_complete/word_0/ca
      -- 
    ca_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_107_store_0_ack_1, ack => testConfigure_CP_0_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	249 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Sample/word_access_start/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Sample/word_access_start/word_0/rr
      -- 
    rr_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(23), ack => ptr_deref_124_load_0_req_0); -- 
    testConfigure_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(30) & testConfigure_CP_0_elements(249);
      gj_testConfigure_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Sample/word_access_start/$exit
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Sample/word_access_start/word_0/ra
      -- 
    ra_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_124_load_0_ack_0, ack => testConfigure_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	249 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	31 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/word_access_complete/$exit
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/ptr_deref_124_Merge/$entry
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/ptr_deref_124_Merge/$exit
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/ptr_deref_124_Merge/merge_req
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/ptr_deref_124_Merge/merge_ack
      -- 
    ca_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_124_load_0_ack_1, ack => testConfigure_CP_0_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	249 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_update_start_
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_Update/cr
      -- 
    ra_407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_132_inst_ack_0, ack => testConfigure_CP_0_elements(26)); -- 
    cr_411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(26), ack => RPIPE_ConvTranspose_input_pipe_132_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_Sample/rr
      -- 
    ca_412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_132_inst_ack_1, ack => testConfigure_CP_0_elements(27)); -- 
    rr_420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(27), ack => type_cast_136_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_Sample/ra
      -- 
    ra_421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_136_inst_ack_0, ack => testConfigure_CP_0_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	249 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_Update/ca
      -- 
    ca_426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_136_inst_ack_1, ack => testConfigure_CP_0_elements(29)); -- 
    -- CP-element group 30:  transition  delay-element  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	21 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	23 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_ptr_deref_124_delay
      -- 
    -- Element group testConfigure_CP_0_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(21), ack => testConfigure_CP_0_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  branch  join  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	17 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	25 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (10) 
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137__exit__
      -- CP-element group 31: 	 branch_block_stmt_34/if_stmt_138__entry__
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/$exit
      -- CP-element group 31: 	 branch_block_stmt_34/if_stmt_138_dead_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_34/if_stmt_138_eval_test/$entry
      -- CP-element group 31: 	 branch_block_stmt_34/if_stmt_138_eval_test/$exit
      -- CP-element group 31: 	 branch_block_stmt_34/if_stmt_138_eval_test/branch_req
      -- CP-element group 31: 	 branch_block_stmt_34/R_cmp_139_place
      -- CP-element group 31: 	 branch_block_stmt_34/if_stmt_138_if_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_34/if_stmt_138_else_link/$entry
      -- 
    branch_req_435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(31), ack => if_stmt_138_branch_req_0); -- 
    testConfigure_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(29) & testConfigure_CP_0_elements(16) & testConfigure_CP_0_elements(17) & testConfigure_CP_0_elements(22) & testConfigure_CP_0_elements(25);
      gj_testConfigure_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  place  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	234 
    -- CP-element group 32: 	235 
    -- CP-element group 32: 	237 
    -- CP-element group 32: 	238 
    -- CP-element group 32:  members (20) 
      -- CP-element group 32: 	 branch_block_stmt_34/if_stmt_138_if_link/$exit
      -- CP-element group 32: 	 branch_block_stmt_34/if_stmt_138_if_link/if_choice_transition
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/Update/cr
      -- 
    if_choice_transition_440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_138_branch_ack_1, ack => testConfigure_CP_0_elements(32)); -- 
    rr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_78_inst_req_0); -- 
    cr_2668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_78_inst_req_1); -- 
    rr_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_85_inst_req_0); -- 
    cr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_85_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	250 
    -- CP-element group 33: 	251 
    -- CP-element group 33:  members (12) 
      -- CP-element group 33: 	 branch_block_stmt_34/if_stmt_138_else_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_34/if_stmt_138_else_link/else_choice_transition
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/Update/cr
      -- 
    else_choice_transition_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_138_branch_ack_0, ack => testConfigure_CP_0_elements(33)); -- 
    rr_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_148_inst_req_0); -- 
    cr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_148_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	261 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/word_access_start/$exit
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/word_access_start/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/word_access_start/word_0/ra
      -- 
    ra_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_166_store_0_ack_0, ack => testConfigure_CP_0_elements(34)); -- 
    -- CP-element group 35:  branch  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	261 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (15) 
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174__exit__
      -- CP-element group 35: 	 branch_block_stmt_34/if_stmt_175__entry__
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/$exit
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Update/word_access_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Update/word_access_complete/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Update/word_access_complete/word_0/ca
      -- CP-element group 35: 	 branch_block_stmt_34/if_stmt_175_dead_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_34/if_stmt_175_eval_test/$entry
      -- CP-element group 35: 	 branch_block_stmt_34/if_stmt_175_eval_test/$exit
      -- CP-element group 35: 	 branch_block_stmt_34/if_stmt_175_eval_test/branch_req
      -- CP-element group 35: 	 branch_block_stmt_34/R_cmp12223_176_place
      -- CP-element group 35: 	 branch_block_stmt_34/if_stmt_175_if_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_34/if_stmt_175_else_link/$entry
      -- 
    ca_499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_166_store_0_ack_1, ack => testConfigure_CP_0_elements(35)); -- 
    branch_req_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => if_stmt_175_branch_req_0); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	268 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_34/if_stmt_175_if_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_34/if_stmt_175_if_link/if_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_34/forx_xend_bbx_xnph221
      -- CP-element group 36: 	 branch_block_stmt_34/forx_xend_bbx_xnph221_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_34/forx_xend_bbx_xnph221_PhiReq/$exit
      -- 
    if_choice_transition_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_175_branch_ack_1, ack => testConfigure_CP_0_elements(36)); -- 
    -- CP-element group 37:  merge  transition  place  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	265 
    -- CP-element group 37:  members (14) 
      -- CP-element group 37: 	 branch_block_stmt_34/merge_stmt_181__exit__
      -- CP-element group 37: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14
      -- CP-element group 37: 	 branch_block_stmt_34/if_stmt_175_else_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_34/if_stmt_175_else_link/else_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_34/forx_xend_forx_xbody14x_xpreheader
      -- CP-element group 37: 	 branch_block_stmt_34/forx_xend_forx_xbody14x_xpreheader_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_34/forx_xend_forx_xbody14x_xpreheader_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_34/merge_stmt_181_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_34/merge_stmt_181_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_34/merge_stmt_181_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_34/merge_stmt_181_PhiAck/dummy
      -- CP-element group 37: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_184/$entry
      -- CP-element group 37: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/$entry
      -- 
    else_choice_transition_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_175_branch_ack_0, ack => testConfigure_CP_0_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	267 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_Sample/ra
      -- 
    ra_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_200_inst_ack_0, ack => testConfigure_CP_0_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	267 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_Update/ca
      -- 
    ca_535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_200_inst_ack_1, ack => testConfigure_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	267 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	55 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_sample_complete
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_Sample/ack
      -- 
    ack_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_206_index_offset_ack_0, ack => testConfigure_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	267 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (11) 
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_offset_calculated
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_request/$entry
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_request/req
      -- 
    ack_566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_206_index_offset_ack_1, ack => testConfigure_CP_0_elements(41)); -- 
    req_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(41), ack => addr_of_207_final_reg_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_request/$exit
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_request/ack
      -- 
    ack_576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_207_final_reg_ack_0, ack => testConfigure_CP_0_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	267 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	48 
    -- CP-element group 43:  members (19) 
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_complete/ack
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_word_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_address_resized
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_addr_resize/$entry
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_addr_resize/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_addr_resize/base_resize_req
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_addr_resize/base_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_word_addrgen/$entry
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_word_addrgen/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_word_addrgen/root_register_req
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_word_addrgen/root_register_ack
      -- 
    ack_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_207_final_reg_ack_1, ack => testConfigure_CP_0_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	267 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_update_start_
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_Update/cr
      -- 
    ra_590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_210_inst_ack_0, ack => testConfigure_CP_0_elements(44)); -- 
    cr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(44), ack => RPIPE_ConvTranspose_input_pipe_210_inst_req_1); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_Sample/rr
      -- 
    ca_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_210_inst_ack_1, ack => testConfigure_CP_0_elements(45)); -- 
    rr_603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(45), ack => type_cast_214_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_Sample/ra
      -- 
    ra_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_0, ack => testConfigure_CP_0_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	267 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_Update/ca
      -- 
    ca_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_1, ack => testConfigure_CP_0_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	43 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/ptr_deref_217_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/ptr_deref_217_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/ptr_deref_217_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/ptr_deref_217_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/word_access_start/word_0/rr
      -- 
    rr_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(48), ack => ptr_deref_217_store_0_req_0); -- 
    testConfigure_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(43) & testConfigure_CP_0_elements(47);
      gj_testConfigure_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	54 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Sample/word_access_start/word_0/ra
      -- 
    ra_648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_217_store_0_ack_0, ack => testConfigure_CP_0_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	267 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	55 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Update/word_access_complete/word_0/ca
      -- 
    ca_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_217_store_0_ack_1, ack => testConfigure_CP_0_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: 	267 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Sample/word_access_start/word_0/rr
      -- 
    rr_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => ptr_deref_234_load_0_req_0); -- 
    testConfigure_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(54) & testConfigure_CP_0_elements(267);
      gj_testConfigure_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Sample/word_access_start/word_0/ra
      -- 
    ra_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_234_load_0_ack_0, ack => testConfigure_CP_0_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	267 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/word_access_complete/word_0/ca
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/ptr_deref_234_Merge/$entry
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/ptr_deref_234_Merge/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/ptr_deref_234_Merge/merge_req
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/ptr_deref_234_Merge/merge_ack
      -- 
    ca_704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_234_load_0_ack_1, ack => testConfigure_CP_0_elements(53)); -- 
    -- CP-element group 54:  transition  delay-element  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	49 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_ptr_deref_234_delay
      -- 
    -- Element group testConfigure_CP_0_elements(54) is a control-delay.
    cp_element_54_delay: control_delay_element  generic map(name => " 54_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(49), ack => testConfigure_CP_0_elements(54), clk => clk, reset =>reset);
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: 	40 
    -- CP-element group 55: 	50 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240__exit__
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_241__entry__
      -- CP-element group 55: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/$exit
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_241_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_241_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_241_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_241_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_34/R_cmp12_242_place
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_241_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_241_else_link/$entry
      -- 
    branch_req_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => if_stmt_241_branch_req_0); -- 
    testConfigure_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(39) & testConfigure_CP_0_elements(40) & testConfigure_CP_0_elements(50) & testConfigure_CP_0_elements(53);
      gj_testConfigure_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	262 
    -- CP-element group 56: 	263 
    -- CP-element group 56:  members (12) 
      -- CP-element group 56: 	 branch_block_stmt_34/if_stmt_241_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/if_stmt_241_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/Update/cr
      -- 
    if_choice_transition_723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_241_branch_ack_1, ack => testConfigure_CP_0_elements(56)); -- 
    rr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_187_inst_req_0); -- 
    cr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_187_inst_req_1); -- 
    -- CP-element group 57:  merge  transition  place  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	268 
    -- CP-element group 57:  members (13) 
      -- CP-element group 57: 	 branch_block_stmt_34/merge_stmt_247__exit__
      -- CP-element group 57: 	 branch_block_stmt_34/bbx_xnph221x_xloopexit_bbx_xnph221
      -- CP-element group 57: 	 branch_block_stmt_34/if_stmt_241_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_34/if_stmt_241_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_34/forx_xbody14_bbx_xnph221x_xloopexit
      -- CP-element group 57: 	 branch_block_stmt_34/forx_xbody14_bbx_xnph221x_xloopexit_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_34/forx_xbody14_bbx_xnph221x_xloopexit_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_34/merge_stmt_247_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_34/merge_stmt_247_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_34/merge_stmt_247_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_34/merge_stmt_247_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_34/bbx_xnph221x_xloopexit_bbx_xnph221_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_34/bbx_xnph221x_xloopexit_bbx_xnph221_PhiReq/$exit
      -- 
    else_choice_transition_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_241_branch_ack_0, ack => testConfigure_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	268 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_update_start_
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_Update/cr
      -- 
    ra_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_251_inst_ack_0, ack => testConfigure_CP_0_elements(58)); -- 
    cr_745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(58), ack => RPIPE_ConvTranspose_input_pipe_251_inst_req_1); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_Sample/rr
      -- 
    ca_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_251_inst_ack_1, ack => testConfigure_CP_0_elements(59)); -- 
    rr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(59), ack => type_cast_255_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_Sample/ra
      -- 
    ra_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_0, ack => testConfigure_CP_0_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	268 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	269 
    -- CP-element group 61: 	270 
    -- CP-element group 61: 	271 
    -- CP-element group 61:  members (17) 
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256__exit__
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/$exit
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_259/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/Update/cr
      -- 
    ca_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_1, ack => testConfigure_CP_0_elements(61)); -- 
    rr_2929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(61), ack => type_cast_269_inst_req_0); -- 
    cr_2934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(61), ack => type_cast_269_inst_req_1); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	284 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_request/$exit
      -- CP-element group 62: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_request/ack
      -- CP-element group 62: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_sample_completed_
      -- 
    ack_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_276_final_reg_ack_0, ack => testConfigure_CP_0_elements(62)); -- 
    -- CP-element group 63:  join  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	284 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (28) 
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_complete/ack
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_word_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_root_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_address_resized
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_addr_resize/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_addr_resize/$exit
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_addr_resize/base_resize_req
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_addr_resize/base_resize_ack
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_plus_offset/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_plus_offset/$exit
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_plus_offset/sum_rename_req
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_base_plus_offset/sum_rename_ack
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_word_addrgen/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_word_addrgen/$exit
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_word_addrgen/root_register_req
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_word_addrgen/root_register_ack
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/ptr_deref_279_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/ptr_deref_279_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/ptr_deref_279_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/ptr_deref_279_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/word_access_start/word_0/rr
      -- 
    ack_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_276_final_reg_ack_1, ack => testConfigure_CP_0_elements(63)); -- 
    rr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(63), ack => ptr_deref_279_store_0_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Sample/word_access_start/word_0/ra
      -- 
    ra_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_279_store_0_ack_0, ack => testConfigure_CP_0_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	284 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	70 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Update/word_access_complete/word_0/ca
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_279_store_0_ack_1, ack => testConfigure_CP_0_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	284 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_update_start_
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_Update/cr
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_283_inst_ack_0, ack => testConfigure_CP_0_elements(66)); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(66), ack => RPIPE_ConvTranspose_input_pipe_283_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_Sample/rr
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_283_inst_ack_1, ack => testConfigure_CP_0_elements(67)); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(67), ack => type_cast_287_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_Sample/ra
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_287_inst_ack_0, ack => testConfigure_CP_0_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	284 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_Update/ca
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_287_inst_ack_1, ack => testConfigure_CP_0_elements(69)); -- 
    -- CP-element group 70:  branch  join  transition  place  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	65 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (10) 
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300__exit__
      -- CP-element group 70: 	 branch_block_stmt_34/if_stmt_301__entry__
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/$exit
      -- CP-element group 70: 	 branch_block_stmt_34/if_stmt_301_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_34/if_stmt_301_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_34/if_stmt_301_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_34/if_stmt_301_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_34/R_exitcond_302_place
      -- CP-element group 70: 	 branch_block_stmt_34/if_stmt_301_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_34/if_stmt_301_else_link/$entry
      -- 
    branch_req_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(70), ack => if_stmt_301_branch_req_0); -- 
    testConfigure_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(65) & testConfigure_CP_0_elements(69);
      gj_testConfigure_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	285 
    -- CP-element group 71: 	286 
    -- CP-element group 71:  members (12) 
      -- CP-element group 71: 	 branch_block_stmt_34/if_stmt_301_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/if_stmt_301_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/Update/cr
      -- 
    if_choice_transition_893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_301_branch_ack_1, ack => testConfigure_CP_0_elements(71)); -- 
    rr_3014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_311_inst_req_0); -- 
    cr_3019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_311_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	274 
    -- CP-element group 72: 	275 
    -- CP-element group 72: 	277 
    -- CP-element group 72: 	278 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_34/if_stmt_301_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_34/if_stmt_301_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/Update/cr
      -- 
    else_choice_transition_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_301_branch_ack_0, ack => testConfigure_CP_0_elements(72)); -- 
    rr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_265_inst_req_0); -- 
    cr_2960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_265_inst_req_1); -- 
    rr_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_271_inst_req_0); -- 
    cr_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_271_inst_req_1); -- 
    -- CP-element group 73:  join  fork  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	288 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	76 
    -- CP-element group 73: 	79 
    -- CP-element group 73: 	80 
    -- CP-element group 73: 	82 
    -- CP-element group 73: 	86 
    -- CP-element group 73: 	87 
    -- CP-element group 73: 	89 
    -- CP-element group 73: 	93 
    -- CP-element group 73: 	94 
    -- CP-element group 73: 	96 
    -- CP-element group 73: 	97 
    -- CP-element group 73: 	98 
    -- CP-element group 73: 	99 
    -- CP-element group 73: 	100 
    -- CP-element group 73: 	101 
    -- CP-element group 73: 	102 
    -- CP-element group 73: 	105 
    -- CP-element group 73: 	106 
    -- CP-element group 73: 	107 
    -- CP-element group 73: 	108 
    -- CP-element group 73: 	109 
    -- CP-element group 73: 	110 
    -- CP-element group 73: 	111 
    -- CP-element group 73: 	112 
    -- CP-element group 73: 	113 
    -- CP-element group 73: 	116 
    -- CP-element group 73:  members (280) 
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/STORE_padding_313_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/STORE_padding_313_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/STORE_padding_313_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/STORE_padding_313_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Update/word_access_complete/word_0/cr
      -- 
    cr_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => STORE_padding_313_store_0_req_1); -- 
    rr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => STORE_padding_313_store_0_req_0); -- 
    rr_943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => RPIPE_ConvTranspose_input_pipe_317_inst_req_0); -- 
    cr_962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_321_inst_req_1); -- 
    cr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_332_store_0_req_1); -- 
    cr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_340_inst_req_1); -- 
    cr_1090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_351_store_0_req_1); -- 
    cr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_359_inst_req_1); -- 
    cr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_370_store_0_req_1); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_383_load_0_req_1); -- 
    rr_1202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_383_load_0_req_0); -- 
    cr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_395_load_0_req_1); -- 
    rr_1252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_395_load_0_req_0); -- 
    cr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_407_load_0_req_1); -- 
    rr_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_407_load_0_req_0); -- 
    cr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_421_inst_req_1); -- 
    cr_1377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_433_load_0_req_1); -- 
    rr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_433_load_0_req_0); -- 
    cr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_445_load_0_req_1); -- 
    rr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_445_load_0_req_0); -- 
    cr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_457_load_0_req_1); -- 
    rr_1466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_457_load_0_req_0); -- 
    cr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_469_load_0_req_1); -- 
    rr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_469_load_0_req_0); -- 
    cr_1546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_488_inst_req_1); -- 
    testConfigure_CP_0_elements(73) <= testConfigure_CP_0_elements(288);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Sample/word_access_start/word_0/ra
      -- 
    ra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_313_store_0_ack_0, ack => testConfigure_CP_0_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	119 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/STORE_padding_313_Update/word_access_complete/word_0/ca
      -- 
    ca_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_313_store_0_ack_1, ack => testConfigure_CP_0_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	73 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_update_start_
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_Update/cr
      -- 
    ra_944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_317_inst_ack_0, ack => testConfigure_CP_0_elements(76)); -- 
    cr_948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => RPIPE_ConvTranspose_input_pipe_317_inst_req_1); -- 
    -- CP-element group 77:  fork  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	83 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_317_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_Sample/rr
      -- 
    ca_949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_317_inst_ack_1, ack => testConfigure_CP_0_elements(77)); -- 
    rr_957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_321_inst_req_0); -- 
    rr_1021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => RPIPE_ConvTranspose_input_pipe_336_inst_req_0); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_Sample/ra
      -- 
    ra_958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_321_inst_ack_0, ack => testConfigure_CP_0_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	73 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_321_Update/ca
      -- 
    ca_963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_321_inst_ack_1, ack => testConfigure_CP_0_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	73 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/ptr_deref_332_Split/$entry
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/ptr_deref_332_Split/$exit
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/ptr_deref_332_Split/split_req
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/ptr_deref_332_Split/split_ack
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/word_access_start/word_0/rr
      -- 
    rr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(80), ack => ptr_deref_332_store_0_req_0); -- 
    testConfigure_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(79);
      gj_testConfigure_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	117 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/word_access_start/$exit
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/word_access_start/word_0/$exit
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Sample/word_access_start/word_0/ra
      -- 
    ra_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_332_store_0_ack_0, ack => testConfigure_CP_0_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	73 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	119 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Update/word_access_complete/$exit
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Update/word_access_complete/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_Update/word_access_complete/word_0/ca
      -- 
    ca_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_332_store_0_ack_1, ack => testConfigure_CP_0_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_update_start_
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_Update/cr
      -- 
    ra_1022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_336_inst_ack_0, ack => testConfigure_CP_0_elements(83)); -- 
    cr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(83), ack => RPIPE_ConvTranspose_input_pipe_336_inst_req_1); -- 
    -- CP-element group 84:  fork  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	90 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_336_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_Sample/rr
      -- 
    ca_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_336_inst_ack_1, ack => testConfigure_CP_0_elements(84)); -- 
    rr_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => type_cast_340_inst_req_0); -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => RPIPE_ConvTranspose_input_pipe_355_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_Sample/ra
      -- 
    ra_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_340_inst_ack_0, ack => testConfigure_CP_0_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	73 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_340_Update/ca
      -- 
    ca_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_340_inst_ack_1, ack => testConfigure_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	73 
    -- CP-element group 87: 	86 
    -- CP-element group 87: 	117 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/ptr_deref_351_Split/$entry
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/ptr_deref_351_Split/$exit
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/ptr_deref_351_Split/split_req
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/ptr_deref_351_Split/split_ack
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/word_access_start/$entry
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/word_access_start/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/word_access_start/word_0/rr
      -- 
    rr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(87), ack => ptr_deref_351_store_0_req_0); -- 
    testConfigure_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(86) & testConfigure_CP_0_elements(117);
      gj_testConfigure_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	118 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/word_access_start/$exit
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/word_access_start/word_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Sample/word_access_start/word_0/ra
      -- 
    ra_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_351_store_0_ack_0, ack => testConfigure_CP_0_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	73 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	119 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Update/word_access_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Update/word_access_complete/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_Update/word_access_complete/word_0/ca
      -- 
    ca_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_351_store_0_ack_1, ack => testConfigure_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	84 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_update_start_
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_Update/cr
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_355_inst_ack_0, ack => testConfigure_CP_0_elements(90)); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(90), ack => RPIPE_ConvTranspose_input_pipe_355_inst_req_1); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/RPIPE_ConvTranspose_input_pipe_355_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_sample_start_
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_355_inst_ack_1, ack => testConfigure_CP_0_elements(91)); -- 
    rr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(91), ack => type_cast_359_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_sample_completed_
      -- 
    ra_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_359_inst_ack_0, ack => testConfigure_CP_0_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	73 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_359_Update/$exit
      -- 
    ca_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_359_inst_ack_1, ack => testConfigure_CP_0_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	73 
    -- CP-element group 94: 	93 
    -- CP-element group 94: 	118 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/word_access_start/word_0/rr
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/word_access_start/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/word_access_start/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/ptr_deref_370_Split/split_ack
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/ptr_deref_370_Split/split_req
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/ptr_deref_370_Split/$exit
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/ptr_deref_370_Split/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/$entry
      -- 
    rr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => ptr_deref_370_store_0_req_0); -- 
    testConfigure_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(93) & testConfigure_CP_0_elements(118);
      gj_testConfigure_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/word_access_start/word_0/ra
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/word_access_start/$exit
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Sample/$exit
      -- 
    ra_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_370_store_0_ack_0, ack => testConfigure_CP_0_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	73 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	119 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Update/word_access_complete/word_0/ca
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Update/word_access_complete/word_0/$exit
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Update/word_access_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_370_Update/$exit
      -- 
    ca_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_370_store_0_ack_1, ack => testConfigure_CP_0_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	73 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Sample/word_access_start/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Sample/word_access_start/$exit
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Sample/word_access_start/word_0/ra
      -- 
    ra_1203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_383_load_0_ack_0, ack => testConfigure_CP_0_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	73 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	103 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/ptr_deref_383_Merge/merge_ack
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/ptr_deref_383_Merge/merge_req
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/ptr_deref_383_Merge/$exit
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/ptr_deref_383_Merge/$entry
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/word_access_complete/word_0/ca
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/word_access_complete/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/word_access_complete/$exit
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_383_update_completed_
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_383_load_0_ack_1, ack => testConfigure_CP_0_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	73 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Sample/word_access_start/word_0/ra
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Sample/word_access_start/$exit
      -- 
    ra_1253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_395_load_0_ack_0, ack => testConfigure_CP_0_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	73 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/ptr_deref_395_Merge/$entry
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/word_access_complete/word_0/ca
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/ptr_deref_395_Merge/merge_ack
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/ptr_deref_395_Merge/merge_req
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_395_Update/ptr_deref_395_Merge/$exit
      -- 
    ca_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_395_load_0_ack_1, ack => testConfigure_CP_0_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	73 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Sample/word_access_start/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Sample/$exit
      -- 
    ra_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_407_load_0_ack_0, ack => testConfigure_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	73 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/ptr_deref_407_Merge/merge_req
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/ptr_deref_407_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/ptr_deref_407_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/word_access_complete/word_0/ca
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/word_access_complete/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_407_Update/ptr_deref_407_Merge/merge_ack
      -- 
    ca_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_407_load_0_ack_1, ack => testConfigure_CP_0_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	98 
    -- CP-element group 103: 	100 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_sample_start_
      -- 
    rr_1327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(103), ack => type_cast_421_inst_req_0); -- 
    testConfigure_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(98) & testConfigure_CP_0_elements(100) & testConfigure_CP_0_elements(102);
      gj_testConfigure_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_sample_completed_
      -- 
    ra_1328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_421_inst_ack_0, ack => testConfigure_CP_0_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	73 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	119 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_421_update_completed_
      -- 
    ca_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_421_inst_ack_1, ack => testConfigure_CP_0_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	73 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Sample/word_access_start/word_0/ra
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Sample/word_access_start/word_0/$exit
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Sample/word_access_start/$exit
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Sample/$exit
      -- 
    ra_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_433_load_0_ack_0, ack => testConfigure_CP_0_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	73 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	114 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/ptr_deref_433_Merge/merge_ack
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/ptr_deref_433_Merge/merge_req
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/ptr_deref_433_Merge/$exit
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/ptr_deref_433_Merge/$entry
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/word_access_complete/word_0/ca
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/word_access_complete/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/word_access_complete/$exit
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_433_Update/$exit
      -- 
    ca_1378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_433_load_0_ack_1, ack => testConfigure_CP_0_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	73 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Sample/word_access_start/word_0/ra
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Sample/word_access_start/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Sample/word_access_start/$exit
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Sample/$exit
      -- 
    ra_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_445_load_0_ack_0, ack => testConfigure_CP_0_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	73 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	114 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/ptr_deref_445_Merge/merge_ack
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/ptr_deref_445_Merge/merge_req
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/ptr_deref_445_Merge/$exit
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/ptr_deref_445_Merge/$entry
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/word_access_complete/word_0/ca
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/word_access_complete/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/word_access_complete/$exit
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_445_update_completed_
      -- 
    ca_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_445_load_0_ack_1, ack => testConfigure_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	73 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Sample/word_access_start/word_0/ra
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Sample/word_access_start/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Sample/word_access_start/$exit
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Sample/$exit
      -- 
    ra_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_457_load_0_ack_0, ack => testConfigure_CP_0_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	73 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/word_access_complete/word_0/ca
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/word_access_complete/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/word_access_complete/$exit
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/ptr_deref_457_Merge/merge_ack
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/ptr_deref_457_Merge/merge_req
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/ptr_deref_457_Merge/$exit
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_457_Update/ptr_deref_457_Merge/$entry
      -- 
    ca_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_457_load_0_ack_1, ack => testConfigure_CP_0_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	73 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Sample/word_access_start/word_0/ra
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Sample/word_access_start/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Sample/word_access_start/$exit
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Sample/$exit
      -- 
    ra_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_469_load_0_ack_0, ack => testConfigure_CP_0_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	73 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (9) 
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/word_access_complete/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/ptr_deref_469_Merge/merge_req
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/ptr_deref_469_Merge/$exit
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/ptr_deref_469_Merge/$entry
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/word_access_complete/word_0/ca
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/ptr_deref_469_Merge/merge_ack
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_469_Update/word_access_complete/$exit
      -- 
    ca_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_469_load_0_ack_1, ack => testConfigure_CP_0_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	107 
    -- CP-element group 114: 	109 
    -- CP-element group 114: 	111 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_Sample/$entry
      -- 
    rr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(114), ack => type_cast_488_inst_req_0); -- 
    testConfigure_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(107) & testConfigure_CP_0_elements(109) & testConfigure_CP_0_elements(111) & testConfigure_CP_0_elements(113);
      gj_testConfigure_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_sample_completed_
      -- 
    ra_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_488_inst_ack_0, ack => testConfigure_CP_0_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	73 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/type_cast_488_Update/ca
      -- 
    ca_1547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_488_inst_ack_1, ack => testConfigure_CP_0_elements(116)); -- 
    -- CP-element group 117:  transition  delay-element  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	81 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	87 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_332_ptr_deref_351_delay
      -- 
    -- Element group testConfigure_CP_0_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(81), ack => testConfigure_CP_0_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  transition  delay-element  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	94 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/ptr_deref_351_ptr_deref_370_delay
      -- 
    -- Element group testConfigure_CP_0_elements(118) is a control-delay.
    cp_element_118_delay: control_delay_element  generic map(name => " 118_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(88), ack => testConfigure_CP_0_elements(118), clk => clk, reset =>reset);
    -- CP-element group 119:  branch  join  transition  place  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	75 
    -- CP-element group 119: 	82 
    -- CP-element group 119: 	89 
    -- CP-element group 119: 	96 
    -- CP-element group 119: 	105 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (10) 
      -- CP-element group 119: 	 branch_block_stmt_34/if_stmt_502_if_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/if_stmt_502_else_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/if_stmt_502_dead_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/if_stmt_502_eval_test/$entry
      -- CP-element group 119: 	 branch_block_stmt_34/if_stmt_502_eval_test/$exit
      -- CP-element group 119: 	 branch_block_stmt_34/if_stmt_502_eval_test/branch_req
      -- CP-element group 119: 	 branch_block_stmt_34/R_cmp65213_503_place
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501__exit__
      -- CP-element group 119: 	 branch_block_stmt_34/if_stmt_502__entry__
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501/$exit
      -- 
    branch_req_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => if_stmt_502_branch_req_0); -- 
    testConfigure_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(75) & testConfigure_CP_0_elements(82) & testConfigure_CP_0_elements(89) & testConfigure_CP_0_elements(96) & testConfigure_CP_0_elements(105) & testConfigure_CP_0_elements(116);
      gj_testConfigure_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	289 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_502_if_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_502_if_link/if_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_34/forx_xend37_forx_xcond119x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_34/forx_xend37_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_34/forx_xend37_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_502_branch_ack_1, ack => testConfigure_CP_0_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	124 
    -- CP-element group 121: 	125 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_34/if_stmt_502_else_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_34/if_stmt_502_else_link/else_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_529__exit__
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562__entry__
      -- CP-element group 121: 	 branch_block_stmt_34/forx_xend37_bbx_xnph215
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_update_start_
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_34/forx_xend37_bbx_xnph215_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/forx_xend37_bbx_xnph215_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_529_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_529_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_529_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_529_PhiAck/dummy
      -- 
    else_choice_transition_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_502_branch_ack_0, ack => testConfigure_CP_0_elements(121)); -- 
    rr_1601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_542_inst_req_0); -- 
    cr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_542_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	289 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	302 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_34/if_stmt_523_if_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_34/if_stmt_523_if_link/if_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_34/forx_xcond119x_xpreheader_forx_xend180
      -- CP-element group 122: 	 branch_block_stmt_34/forx_xcond119x_xpreheader_forx_xend180_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_34/forx_xcond119x_xpreheader_forx_xend180_PhiReq/$exit
      -- 
    if_choice_transition_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_523_branch_ack_1, ack => testConfigure_CP_0_elements(122)); -- 
    -- CP-element group 123:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	289 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	168 
    -- CP-element group 123: 	169 
    -- CP-element group 123:  members (18) 
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_734__exit__
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772__entry__
      -- CP-element group 123: 	 branch_block_stmt_34/if_stmt_523_else_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_34/if_stmt_523_else_link/else_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_34/forx_xcond119x_xpreheader_bbx_xnph210
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_update_start_
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_34/forx_xcond119x_xpreheader_bbx_xnph210_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/forx_xcond119x_xpreheader_bbx_xnph210_PhiReq/$exit
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_734_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_734_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_734_PhiAck/$exit
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_734_PhiAck/dummy
      -- 
    else_choice_transition_1588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_523_branch_ack_0, ack => testConfigure_CP_0_elements(123)); -- 
    rr_1960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_752_inst_req_0); -- 
    cr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_752_inst_req_1); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_Sample/ra
      -- 
    ra_1602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_542_inst_ack_0, ack => testConfigure_CP_0_elements(124)); -- 
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	121 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	290 
    -- CP-element group 125:  members (9) 
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562__exit__
      -- CP-element group 125: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/$exit
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_534_to_assign_stmt_562/type_cast_542_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67_PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_565/$entry
      -- CP-element group 125: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/$entry
      -- 
    ca_1607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_542_inst_ack_1, ack => testConfigure_CP_0_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	295 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	165 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_sample_complete
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_Sample/ack
      -- 
    ack_1636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_577_index_offset_ack_0, ack => testConfigure_CP_0_elements(126)); -- 
    -- CP-element group 127:  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	295 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (11) 
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_root_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_offset_calculated
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_Update/ack
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_base_plus_offset/$entry
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_base_plus_offset/$exit
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_base_plus_offset/sum_rename_req
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_base_plus_offset/sum_rename_ack
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_request/$entry
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_request/req
      -- 
    ack_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_577_index_offset_ack_1, ack => testConfigure_CP_0_elements(127)); -- 
    req_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(127), ack => addr_of_578_final_reg_req_0); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_request/$exit
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_request/ack
      -- 
    ack_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_578_final_reg_ack_0, ack => testConfigure_CP_0_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	295 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	162 
    -- CP-element group 129:  members (19) 
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_complete/ack
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_word_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_root_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_address_resized
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_addr_resize/$entry
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_addr_resize/$exit
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_addr_resize/base_resize_req
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_addr_resize/base_resize_ack
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_plus_offset/$entry
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_plus_offset/$exit
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_plus_offset/sum_rename_req
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_base_plus_offset/sum_rename_ack
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_word_addrgen/$entry
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_word_addrgen/$exit
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_word_addrgen/root_register_req
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_word_addrgen/root_register_ack
      -- 
    ack_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_578_final_reg_ack_1, ack => testConfigure_CP_0_elements(129)); -- 
    -- CP-element group 130:  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	295 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_update_start_
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_Sample/ra
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_Update/cr
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_581_inst_ack_0, ack => testConfigure_CP_0_elements(130)); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(130), ack => RPIPE_ConvTranspose_input_pipe_581_inst_req_1); -- 
    -- CP-element group 131:  fork  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (9) 
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_Sample/rr
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_581_inst_ack_1, ack => testConfigure_CP_0_elements(131)); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => type_cast_585_inst_req_0); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => RPIPE_ConvTranspose_input_pipe_594_inst_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_0, ack => testConfigure_CP_0_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	295 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	162 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_Update/ca
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_1, ack => testConfigure_CP_0_elements(133)); -- 
    -- CP-element group 134:  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_update_start_
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_Update/cr
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_594_inst_ack_0, ack => testConfigure_CP_0_elements(134)); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(134), ack => RPIPE_ConvTranspose_input_pipe_594_inst_req_1); -- 
    -- CP-element group 135:  fork  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (9) 
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_594_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_Sample/rr
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_Sample/rr
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_594_inst_ack_1, ack => testConfigure_CP_0_elements(135)); -- 
    rr_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => type_cast_598_inst_req_0); -- 
    rr_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => RPIPE_ConvTranspose_input_pipe_612_inst_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_Sample/ra
      -- 
    ra_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_0, ack => testConfigure_CP_0_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	295 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	162 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_Update/ca
      -- 
    ca_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_1, ack => testConfigure_CP_0_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_update_start_
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_Update/cr
      -- 
    ra_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_612_inst_ack_0, ack => testConfigure_CP_0_elements(138)); -- 
    cr_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(138), ack => RPIPE_ConvTranspose_input_pipe_612_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	142 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_612_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_Sample/rr
      -- 
    ca_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_612_inst_ack_1, ack => testConfigure_CP_0_elements(139)); -- 
    rr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => type_cast_616_inst_req_0); -- 
    rr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => RPIPE_ConvTranspose_input_pipe_630_inst_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_Sample/ra
      -- 
    ra_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_0, ack => testConfigure_CP_0_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	295 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	162 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_Update/ca
      -- 
    ca_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_1, ack => testConfigure_CP_0_elements(141)); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_update_start_
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_Update/cr
      -- 
    ra_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_630_inst_ack_0, ack => testConfigure_CP_0_elements(142)); -- 
    cr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(142), ack => RPIPE_ConvTranspose_input_pipe_630_inst_req_1); -- 
    -- CP-element group 143:  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: 	146 
    -- CP-element group 143:  members (9) 
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_630_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_Sample/rr
      -- 
    ca_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_630_inst_ack_1, ack => testConfigure_CP_0_elements(143)); -- 
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => type_cast_634_inst_req_0); -- 
    rr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => RPIPE_ConvTranspose_input_pipe_648_inst_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_Sample/ra
      -- 
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_634_inst_ack_0, ack => testConfigure_CP_0_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	295 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	162 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_Update/ca
      -- 
    ca_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_634_inst_ack_1, ack => testConfigure_CP_0_elements(145)); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	143 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (6) 
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_update_start_
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_Update/cr
      -- 
    ra_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_648_inst_ack_0, ack => testConfigure_CP_0_elements(146)); -- 
    cr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(146), ack => RPIPE_ConvTranspose_input_pipe_648_inst_req_1); -- 
    -- CP-element group 147:  fork  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147: 	150 
    -- CP-element group 147:  members (9) 
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_648_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_Sample/rr
      -- 
    ca_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_648_inst_ack_1, ack => testConfigure_CP_0_elements(147)); -- 
    rr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => type_cast_652_inst_req_0); -- 
    rr_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => RPIPE_ConvTranspose_input_pipe_666_inst_req_0); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_Sample/ra
      -- 
    ra_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_0, ack => testConfigure_CP_0_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	295 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	162 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_Update/ca
      -- 
    ca_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_1, ack => testConfigure_CP_0_elements(149)); -- 
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	147 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_update_start_
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_Update/cr
      -- 
    ra_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_666_inst_ack_0, ack => testConfigure_CP_0_elements(150)); -- 
    cr_1809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(150), ack => RPIPE_ConvTranspose_input_pipe_666_inst_req_1); -- 
    -- CP-element group 151:  fork  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	154 
    -- CP-element group 151:  members (9) 
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_666_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_Sample/rr
      -- 
    ca_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_666_inst_ack_1, ack => testConfigure_CP_0_elements(151)); -- 
    rr_1818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => type_cast_670_inst_req_0); -- 
    rr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => RPIPE_ConvTranspose_input_pipe_684_inst_req_0); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_Sample/ra
      -- 
    ra_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_670_inst_ack_0, ack => testConfigure_CP_0_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	295 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	162 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_Update/ca
      -- 
    ca_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_670_inst_ack_1, ack => testConfigure_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	151 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_update_start_
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_Update/cr
      -- 
    ra_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_684_inst_ack_0, ack => testConfigure_CP_0_elements(154)); -- 
    cr_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(154), ack => RPIPE_ConvTranspose_input_pipe_684_inst_req_1); -- 
    -- CP-element group 155:  fork  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_684_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_Sample/rr
      -- 
    ca_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_684_inst_ack_1, ack => testConfigure_CP_0_elements(155)); -- 
    rr_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => type_cast_688_inst_req_0); -- 
    rr_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => RPIPE_ConvTranspose_input_pipe_702_inst_req_0); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_Sample/ra
      -- 
    ra_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_0, ack => testConfigure_CP_0_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	295 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_Update/ca
      -- 
    ca_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_1, ack => testConfigure_CP_0_elements(157)); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_update_start_
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_Update/cr
      -- 
    ra_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_702_inst_ack_0, ack => testConfigure_CP_0_elements(158)); -- 
    cr_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(158), ack => RPIPE_ConvTranspose_input_pipe_702_inst_req_1); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_702_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_Sample/rr
      -- 
    ca_1866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_702_inst_ack_1, ack => testConfigure_CP_0_elements(159)); -- 
    rr_1874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(159), ack => type_cast_706_inst_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_Sample/ra
      -- 
    ra_1875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_706_inst_ack_0, ack => testConfigure_CP_0_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	295 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_Update/ca
      -- 
    ca_1880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_706_inst_ack_1, ack => testConfigure_CP_0_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	129 
    -- CP-element group 162: 	133 
    -- CP-element group 162: 	137 
    -- CP-element group 162: 	141 
    -- CP-element group 162: 	145 
    -- CP-element group 162: 	149 
    -- CP-element group 162: 	153 
    -- CP-element group 162: 	157 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (9) 
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/ptr_deref_714_Split/$entry
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/ptr_deref_714_Split/$exit
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/ptr_deref_714_Split/split_req
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/ptr_deref_714_Split/split_ack
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/word_access_start/$entry
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/word_access_start/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/word_access_start/word_0/rr
      -- 
    rr_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(162), ack => ptr_deref_714_store_0_req_0); -- 
    testConfigure_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(129) & testConfigure_CP_0_elements(133) & testConfigure_CP_0_elements(137) & testConfigure_CP_0_elements(141) & testConfigure_CP_0_elements(145) & testConfigure_CP_0_elements(149) & testConfigure_CP_0_elements(153) & testConfigure_CP_0_elements(157) & testConfigure_CP_0_elements(161);
      gj_testConfigure_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/word_access_start/$exit
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/word_access_start/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Sample/word_access_start/word_0/ra
      -- 
    ra_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_714_store_0_ack_0, ack => testConfigure_CP_0_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	295 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Update/word_access_complete/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Update/word_access_complete/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Update/word_access_complete/word_0/ca
      -- 
    ca_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_714_store_0_ack_1, ack => testConfigure_CP_0_elements(164)); -- 
    -- CP-element group 165:  branch  join  transition  place  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	126 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (10) 
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727__exit__
      -- CP-element group 165: 	 branch_block_stmt_34/if_stmt_728__entry__
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/$exit
      -- CP-element group 165: 	 branch_block_stmt_34/if_stmt_728_dead_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_34/if_stmt_728_eval_test/$entry
      -- CP-element group 165: 	 branch_block_stmt_34/if_stmt_728_eval_test/$exit
      -- CP-element group 165: 	 branch_block_stmt_34/if_stmt_728_eval_test/branch_req
      -- CP-element group 165: 	 branch_block_stmt_34/R_exitcond10_729_place
      -- CP-element group 165: 	 branch_block_stmt_34/if_stmt_728_if_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_34/if_stmt_728_else_link/$entry
      -- 
    branch_req_1938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(165), ack => if_stmt_728_branch_req_0); -- 
    testConfigure_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(126) & testConfigure_CP_0_elements(164);
      gj_testConfigure_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  merge  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	289 
    -- CP-element group 166:  members (13) 
      -- CP-element group 166: 	 branch_block_stmt_34/merge_stmt_508__exit__
      -- CP-element group 166: 	 branch_block_stmt_34/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_728_if_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_728_if_link/if_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_34/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit
      -- CP-element group 166: 	 branch_block_stmt_34/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_34/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 166: 	 branch_block_stmt_34/merge_stmt_508_PhiReqMerge
      -- CP-element group 166: 	 branch_block_stmt_34/merge_stmt_508_PhiAck/$entry
      -- CP-element group 166: 	 branch_block_stmt_34/merge_stmt_508_PhiAck/$exit
      -- CP-element group 166: 	 branch_block_stmt_34/merge_stmt_508_PhiAck/dummy
      -- CP-element group 166: 	 branch_block_stmt_34/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_34/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_728_branch_ack_1, ack => testConfigure_CP_0_elements(166)); -- 
    -- CP-element group 167:  fork  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	291 
    -- CP-element group 167: 	292 
    -- CP-element group 167:  members (12) 
      -- CP-element group 167: 	 branch_block_stmt_34/if_stmt_728_else_link/$exit
      -- CP-element group 167: 	 branch_block_stmt_34/if_stmt_728_else_link/else_choice_transition
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_728_branch_ack_0, ack => testConfigure_CP_0_elements(167)); -- 
    rr_3091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_571_inst_req_0); -- 
    cr_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_571_inst_req_1); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	123 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_Sample/ra
      -- 
    ra_1961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_752_inst_ack_0, ack => testConfigure_CP_0_elements(168)); -- 
    -- CP-element group 169:  transition  place  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	123 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	296 
    -- CP-element group 169:  members (9) 
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772__exit__
      -- CP-element group 169: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/$exit
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_739_to_assign_stmt_772/type_cast_752_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126_PhiReq/$entry
      -- CP-element group 169: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_775/$entry
      -- CP-element group 169: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/$entry
      -- 
    ca_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_752_inst_ack_1, ack => testConfigure_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	301 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	209 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_sample_complete
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_Sample/ack
      -- 
    ack_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_787_index_offset_ack_0, ack => testConfigure_CP_0_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	301 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (11) 
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_root_address_calculated
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_offset_calculated
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_Update/ack
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_base_plus_offset/$entry
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_base_plus_offset/$exit
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_base_plus_offset/sum_rename_req
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_base_plus_offset/sum_rename_ack
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_request/$entry
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_request/req
      -- 
    ack_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_787_index_offset_ack_1, ack => testConfigure_CP_0_elements(171)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(171), ack => addr_of_788_final_reg_req_0); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_request/$exit
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_request/ack
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_788_final_reg_ack_0, ack => testConfigure_CP_0_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	301 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	206 
    -- CP-element group 173:  members (19) 
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_plus_offset/$exit
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_root_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_addr_resize/$entry
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_addr_resize/$exit
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_address_resized
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_addr_resize/base_resize_req
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_addr_resize/base_resize_ack
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_word_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_plus_offset/$entry
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_word_addrgen/root_register_ack
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_word_addrgen/root_register_req
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_word_addrgen/$exit
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_word_addrgen/$entry
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_plus_offset/sum_rename_ack
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_base_plus_offset/sum_rename_req
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_complete/$exit
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_complete/ack
      -- 
    ack_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_788_final_reg_ack_1, ack => testConfigure_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	301 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (6) 
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_update_start_
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_Sample/ra
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_Update/cr
      -- 
    ra_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_791_inst_ack_0, ack => testConfigure_CP_0_elements(174)); -- 
    cr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(174), ack => RPIPE_ConvTranspose_input_pipe_791_inst_req_1); -- 
    -- CP-element group 175:  fork  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: 	178 
    -- CP-element group 175:  members (9) 
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_Sample/rr
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_Sample/rr
      -- 
    ca_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_791_inst_ack_1, ack => testConfigure_CP_0_elements(175)); -- 
    rr_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => type_cast_795_inst_req_0); -- 
    rr_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => RPIPE_ConvTranspose_input_pipe_804_inst_req_0); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_Sample/ra
      -- 
    ra_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_795_inst_ack_0, ack => testConfigure_CP_0_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	301 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	206 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_Update/ca
      -- 
    ca_2043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_795_inst_ack_1, ack => testConfigure_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	175 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (6) 
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_update_start_
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_Sample/ra
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_Update/cr
      -- 
    ra_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_804_inst_ack_0, ack => testConfigure_CP_0_elements(178)); -- 
    cr_2056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(178), ack => RPIPE_ConvTranspose_input_pipe_804_inst_req_1); -- 
    -- CP-element group 179:  fork  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: 	182 
    -- CP-element group 179:  members (9) 
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_804_Update/ca
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_Sample/rr
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_Sample/rr
      -- 
    ca_2057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_804_inst_ack_1, ack => testConfigure_CP_0_elements(179)); -- 
    rr_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => type_cast_808_inst_req_0); -- 
    rr_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => RPIPE_ConvTranspose_input_pipe_822_inst_req_0); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_Sample/ra
      -- 
    ra_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_808_inst_ack_0, ack => testConfigure_CP_0_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	301 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	206 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_Update/ca
      -- 
    ca_2071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_808_inst_ack_1, ack => testConfigure_CP_0_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	179 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (6) 
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_update_start_
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_Sample/ra
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_Update/cr
      -- 
    ra_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_822_inst_ack_0, ack => testConfigure_CP_0_elements(182)); -- 
    cr_2084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(182), ack => RPIPE_ConvTranspose_input_pipe_822_inst_req_1); -- 
    -- CP-element group 183:  fork  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183: 	186 
    -- CP-element group 183:  members (9) 
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_822_Update/ca
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_Sample/rr
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_Sample/rr
      -- 
    ca_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_822_inst_ack_1, ack => testConfigure_CP_0_elements(183)); -- 
    rr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => type_cast_826_inst_req_0); -- 
    rr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => RPIPE_ConvTranspose_input_pipe_840_inst_req_0); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_Sample/ra
      -- 
    ra_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_826_inst_ack_0, ack => testConfigure_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	301 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	206 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_Update/ca
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_826_inst_ack_1, ack => testConfigure_CP_0_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	183 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_update_start_
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_Update/cr
      -- 
    ra_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_840_inst_ack_0, ack => testConfigure_CP_0_elements(186)); -- 
    cr_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(186), ack => RPIPE_ConvTranspose_input_pipe_840_inst_req_1); -- 
    -- CP-element group 187:  fork  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	190 
    -- CP-element group 187:  members (9) 
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_840_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_Sample/rr
      -- 
    ca_2113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_840_inst_ack_1, ack => testConfigure_CP_0_elements(187)); -- 
    rr_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => type_cast_844_inst_req_0); -- 
    rr_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => RPIPE_ConvTranspose_input_pipe_858_inst_req_0); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_Sample/ra
      -- 
    ra_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_844_inst_ack_0, ack => testConfigure_CP_0_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	301 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	206 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_Update/ca
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_update_completed_
      -- 
    ca_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_844_inst_ack_1, ack => testConfigure_CP_0_elements(189)); -- 
    -- CP-element group 190:  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	187 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (6) 
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_Sample/ra
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_update_start_
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_sample_completed_
      -- 
    ra_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_858_inst_ack_0, ack => testConfigure_CP_0_elements(190)); -- 
    cr_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(190), ack => RPIPE_ConvTranspose_input_pipe_858_inst_req_1); -- 
    -- CP-element group 191:  fork  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191: 	194 
    -- CP-element group 191:  members (9) 
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_Sample/rr
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_Update/ca
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_858_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_Sample/rr
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_sample_start_
      -- 
    ca_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_858_inst_ack_1, ack => testConfigure_CP_0_elements(191)); -- 
    rr_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => type_cast_862_inst_req_0); -- 
    rr_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => RPIPE_ConvTranspose_input_pipe_876_inst_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_Sample/ra
      -- 
    ra_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_862_inst_ack_0, ack => testConfigure_CP_0_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	301 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	206 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_Update/ca
      -- 
    ca_2155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_862_inst_ack_1, ack => testConfigure_CP_0_elements(193)); -- 
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	191 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_Update/cr
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_update_start_
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_sample_completed_
      -- 
    ra_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_876_inst_ack_0, ack => testConfigure_CP_0_elements(194)); -- 
    cr_2168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(194), ack => RPIPE_ConvTranspose_input_pipe_876_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195: 	198 
    -- CP-element group 195:  members (9) 
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_876_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_sample_start_
      -- 
    ca_2169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_876_inst_ack_1, ack => testConfigure_CP_0_elements(195)); -- 
    rr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => type_cast_880_inst_req_0); -- 
    rr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => RPIPE_ConvTranspose_input_pipe_894_inst_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_Sample/ra
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_Sample/$exit
      -- 
    ra_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_0, ack => testConfigure_CP_0_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	301 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	206 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_Update/ca
      -- 
    ca_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_1, ack => testConfigure_CP_0_elements(197)); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	195 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_Update/cr
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_update_start_
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_sample_completed_
      -- 
    ra_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_894_inst_ack_0, ack => testConfigure_CP_0_elements(198)); -- 
    cr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(198), ack => RPIPE_ConvTranspose_input_pipe_894_inst_req_1); -- 
    -- CP-element group 199:  fork  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: 	202 
    -- CP-element group 199:  members (9) 
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_894_update_completed_
      -- 
    ca_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_894_inst_ack_1, ack => testConfigure_CP_0_elements(199)); -- 
    rr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => type_cast_898_inst_req_0); -- 
    rr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => RPIPE_ConvTranspose_input_pipe_912_inst_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_sample_completed_
      -- 
    ra_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_0, ack => testConfigure_CP_0_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	301 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	206 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_Update/ca
      -- CP-element group 201: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_update_completed_
      -- 
    ca_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_1, ack => testConfigure_CP_0_elements(201)); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	199 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_update_start_
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_Update/cr
      -- 
    ra_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_912_inst_ack_0, ack => testConfigure_CP_0_elements(202)); -- 
    cr_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(202), ack => RPIPE_ConvTranspose_input_pipe_912_inst_req_1); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_912_Update/ca
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_Sample/rr
      -- 
    ca_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_912_inst_ack_1, ack => testConfigure_CP_0_elements(203)); -- 
    rr_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => type_cast_916_inst_req_0); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_Sample/ra
      -- 
    ra_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_0, ack => testConfigure_CP_0_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	301 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_Update/ca
      -- CP-element group 205: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_Update/$exit
      -- 
    ca_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_1, ack => testConfigure_CP_0_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	173 
    -- CP-element group 206: 	177 
    -- CP-element group 206: 	181 
    -- CP-element group 206: 	185 
    -- CP-element group 206: 	189 
    -- CP-element group 206: 	193 
    -- CP-element group 206: 	197 
    -- CP-element group 206: 	201 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (9) 
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/word_access_start/word_0/rr
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/word_access_start/word_0/$entry
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/word_access_start/$entry
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/ptr_deref_924_Split/split_ack
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/ptr_deref_924_Split/split_req
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/ptr_deref_924_Split/$exit
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/ptr_deref_924_Split/$entry
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/$entry
      -- 
    rr_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(206), ack => ptr_deref_924_store_0_req_0); -- 
    testConfigure_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(173) & testConfigure_CP_0_elements(177) & testConfigure_CP_0_elements(181) & testConfigure_CP_0_elements(185) & testConfigure_CP_0_elements(189) & testConfigure_CP_0_elements(193) & testConfigure_CP_0_elements(197) & testConfigure_CP_0_elements(201) & testConfigure_CP_0_elements(205);
      gj_testConfigure_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/word_access_start/word_0/ra
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/word_access_start/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/word_access_start/$exit
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Sample/$exit
      -- 
    ra_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_924_store_0_ack_0, ack => testConfigure_CP_0_elements(207)); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	301 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Update/word_access_complete/word_0/ca
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Update/word_access_complete/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Update/word_access_complete/$exit
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Update/$exit
      -- 
    ca_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_924_store_0_ack_1, ack => testConfigure_CP_0_elements(208)); -- 
    -- CP-element group 209:  branch  join  transition  place  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	170 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (10) 
      -- CP-element group 209: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937__exit__
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_938__entry__
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_938_else_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_938_if_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_938_eval_test/branch_req
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_938_eval_test/$exit
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_938_eval_test/$entry
      -- CP-element group 209: 	 branch_block_stmt_34/if_stmt_938_dead_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_34/R_exitcond19_939_place
      -- CP-element group 209: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/$exit
      -- 
    branch_req_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(209), ack => if_stmt_938_branch_req_0); -- 
    testConfigure_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(170) & testConfigure_CP_0_elements(208);
      gj_testConfigure_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  merge  transition  place  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	302 
    -- CP-element group 210:  members (13) 
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_944__exit__
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xend180x_xloopexit_forx_xend180
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_938_if_link/if_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_938_if_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xbody126_forx_xend180x_xloopexit
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xbody126_forx_xend180x_xloopexit_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xbody126_forx_xend180x_xloopexit_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_944_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_944_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_944_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_34/merge_stmt_944_PhiAck/dummy
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xend180x_xloopexit_forx_xend180_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/forx_xend180x_xloopexit_forx_xend180_PhiReq/$exit
      -- 
    if_choice_transition_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_938_branch_ack_1, ack => testConfigure_CP_0_elements(210)); -- 
    -- CP-element group 211:  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	297 
    -- CP-element group 211: 	298 
    -- CP-element group 211:  members (12) 
      -- CP-element group 211: 	 branch_block_stmt_34/if_stmt_938_else_link/else_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_34/if_stmt_938_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_938_branch_ack_0, ack => testConfigure_CP_0_elements(211)); -- 
    rr_3145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_781_inst_req_0); -- 
    cr_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_781_inst_req_1); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	303 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (5) 
      -- CP-element group 212: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Sample/word_access_start/$exit
      -- CP-element group 212: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Sample/word_access_start/word_0/ra
      -- CP-element group 212: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Sample/word_access_start/word_0/$exit
      -- CP-element group 212: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_sample_completed_
      -- 
    ra_2345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_957_load_0_ack_0, ack => testConfigure_CP_0_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	303 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	218 
    -- CP-element group 213:  members (9) 
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/word_access_complete/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/word_access_complete/word_0/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/word_access_complete/word_0/ca
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/ptr_deref_957_Merge/$entry
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/ptr_deref_957_Merge/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/ptr_deref_957_Merge/merge_req
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/ptr_deref_957_Merge/merge_ack
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_update_completed_
      -- 
    ca_2356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_957_load_0_ack_1, ack => testConfigure_CP_0_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	303 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (5) 
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Sample/word_access_start/$exit
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Sample/word_access_start/word_0/$exit
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Sample/word_access_start/word_0/ra
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_sample_completed_
      -- 
    ra_2395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_969_load_0_ack_0, ack => testConfigure_CP_0_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	303 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	218 
    -- CP-element group 215:  members (9) 
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/ptr_deref_969_Merge/merge_ack
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/ptr_deref_969_Merge/merge_req
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/ptr_deref_969_Merge/$exit
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/ptr_deref_969_Merge/$entry
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/word_access_complete/word_0/ca
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/word_access_complete/word_0/$exit
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/word_access_complete/$exit
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/$exit
      -- 
    ca_2406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_969_load_0_ack_1, ack => testConfigure_CP_0_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	303 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (5) 
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Sample/word_access_start/word_0/$exit
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Sample/word_access_start/word_0/ra
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Sample/word_access_start/$exit
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_sample_completed_
      -- 
    ra_2445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_981_load_0_ack_0, ack => testConfigure_CP_0_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	303 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (9) 
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/word_access_complete/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/word_access_complete/word_0/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/ptr_deref_981_Merge/merge_ack
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/ptr_deref_981_Merge/merge_req
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/ptr_deref_981_Merge/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/ptr_deref_981_Merge/$entry
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/word_access_complete/word_0/ca
      -- 
    ca_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_981_load_0_ack_1, ack => testConfigure_CP_0_elements(217)); -- 
    -- CP-element group 218:  branch  join  transition  place  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	213 
    -- CP-element group 218: 	215 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (10) 
      -- CP-element group 218: 	 branch_block_stmt_34/if_stmt_999_eval_test/$exit
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998__exit__
      -- CP-element group 218: 	 branch_block_stmt_34/if_stmt_999__entry__
      -- CP-element group 218: 	 branch_block_stmt_34/R_cmp191204_1000_place
      -- CP-element group 218: 	 branch_block_stmt_34/if_stmt_999_eval_test/branch_req
      -- CP-element group 218: 	 branch_block_stmt_34/if_stmt_999_if_link/$entry
      -- CP-element group 218: 	 branch_block_stmt_34/if_stmt_999_else_link/$entry
      -- CP-element group 218: 	 branch_block_stmt_34/if_stmt_999_eval_test/$entry
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/$exit
      -- CP-element group 218: 	 branch_block_stmt_34/if_stmt_999_dead_link/$entry
      -- 
    branch_req_2469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(218), ack => if_stmt_999_branch_req_0); -- 
    testConfigure_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(213) & testConfigure_CP_0_elements(215) & testConfigure_CP_0_elements(217);
      gj_testConfigure_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219: 	222 
    -- CP-element group 219:  members (18) 
      -- CP-element group 219: 	 branch_block_stmt_34/merge_stmt_1005__exit__
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040__entry__
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_Sample/rr
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_999_if_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_999_if_link/if_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_update_start_
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/forx_xend180_bbx_xnph
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_Update/cr
      -- CP-element group 219: 	 branch_block_stmt_34/forx_xend180_bbx_xnph_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/forx_xend180_bbx_xnph_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_34/merge_stmt_1005_PhiReqMerge
      -- CP-element group 219: 	 branch_block_stmt_34/merge_stmt_1005_PhiAck/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/merge_stmt_1005_PhiAck/$exit
      -- CP-element group 219: 	 branch_block_stmt_34/merge_stmt_1005_PhiAck/dummy
      -- 
    if_choice_transition_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_999_branch_ack_1, ack => testConfigure_CP_0_elements(219)); -- 
    rr_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_1026_inst_req_0); -- 
    cr_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_1026_inst_req_1); -- 
    -- CP-element group 220:  transition  place  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	310 
    -- CP-element group 220:  members (5) 
      -- CP-element group 220: 	 branch_block_stmt_34/if_stmt_999_else_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_34/if_stmt_999_else_link/else_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_34/forx_xend180_forx_xend200
      -- CP-element group 220: 	 branch_block_stmt_34/forx_xend180_forx_xend200_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_34/forx_xend180_forx_xend200_PhiReq/$exit
      -- 
    else_choice_transition_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_999_branch_ack_0, ack => testConfigure_CP_0_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_Sample/ra
      -- CP-element group 221: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_sample_completed_
      -- 
    ra_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1026_inst_ack_0, ack => testConfigure_CP_0_elements(221)); -- 
    -- CP-element group 222:  transition  place  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	219 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	304 
    -- CP-element group 222:  members (9) 
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040__exit__
      -- CP-element group 222: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_Update/ca
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/$exit
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_1011_to_assign_stmt_1040/type_cast_1026_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193_PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1043/$entry
      -- CP-element group 222: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/$entry
      -- 
    ca_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1026_inst_ack_1, ack => testConfigure_CP_0_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	309 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	229 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_sample_complete
      -- 
    ack_2526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1055_index_offset_ack_0, ack => testConfigure_CP_0_elements(223)); -- 
    -- CP-element group 224:  transition  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	309 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (11) 
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_base_plus_offset/sum_rename_req
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_base_plus_offset/$exit
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_base_plus_offset/sum_rename_ack
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_base_plus_offset/$entry
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_Update/ack
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_offset_calculated
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_root_address_calculated
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_request/req
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_request/$entry
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_sample_start_
      -- 
    ack_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1055_index_offset_ack_1, ack => testConfigure_CP_0_elements(224)); -- 
    req_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(224), ack => addr_of_1056_final_reg_req_0); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_request/ack
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_request/$exit
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_sample_completed_
      -- 
    ack_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1056_final_reg_ack_0, ack => testConfigure_CP_0_elements(225)); -- 
    -- CP-element group 226:  join  fork  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	309 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (28) 
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_addr_resize/$exit
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_addr_resize/base_resize_req
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_addr_resize/$entry
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_word_addrgen/$entry
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_word_addrgen/$exit
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_plus_offset/sum_rename_ack
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/word_access_start/word_0/rr
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_address_resized
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_complete/ack
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/word_access_start/word_0/$entry
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_root_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_plus_offset/sum_rename_req
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_plus_offset/$exit
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_complete/$exit
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/word_access_start/$entry
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_word_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/ptr_deref_1059_Split/split_ack
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_word_addrgen/root_register_ack
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_plus_offset/$entry
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/ptr_deref_1059_Split/split_req
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/ptr_deref_1059_Split/$exit
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/ptr_deref_1059_Split/$entry
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_word_addrgen/root_register_req
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_base_addr_resize/base_resize_ack
      -- 
    ack_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1056_final_reg_ack_1, ack => testConfigure_CP_0_elements(226)); -- 
    rr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(226), ack => ptr_deref_1059_store_0_req_0); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/word_access_start/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/word_access_start/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Sample/word_access_start/word_0/ra
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_sample_completed_
      -- 
    ra_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1059_store_0_ack_0, ack => testConfigure_CP_0_elements(227)); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	309 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Update/word_access_complete/$exit
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Update/word_access_complete/word_0/$exit
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Update/word_access_complete/word_0/ca
      -- 
    ca_2596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1059_store_0_ack_1, ack => testConfigure_CP_0_elements(228)); -- 
    -- CP-element group 229:  branch  join  transition  place  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	223 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (10) 
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073__exit__
      -- CP-element group 229: 	 branch_block_stmt_34/if_stmt_1074__entry__
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/$exit
      -- CP-element group 229: 	 branch_block_stmt_34/if_stmt_1074_dead_link/$entry
      -- CP-element group 229: 	 branch_block_stmt_34/if_stmt_1074_eval_test/$entry
      -- CP-element group 229: 	 branch_block_stmt_34/if_stmt_1074_eval_test/$exit
      -- CP-element group 229: 	 branch_block_stmt_34/if_stmt_1074_eval_test/branch_req
      -- CP-element group 229: 	 branch_block_stmt_34/R_exitcond20_1075_place
      -- CP-element group 229: 	 branch_block_stmt_34/if_stmt_1074_if_link/$entry
      -- CP-element group 229: 	 branch_block_stmt_34/if_stmt_1074_else_link/$entry
      -- 
    branch_req_2604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => if_stmt_1074_branch_req_0); -- 
    testConfigure_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(223) & testConfigure_CP_0_elements(228);
      gj_testConfigure_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  merge  transition  place  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	310 
    -- CP-element group 230:  members (13) 
      -- CP-element group 230: 	 branch_block_stmt_34/merge_stmt_1080__exit__
      -- CP-element group 230: 	 branch_block_stmt_34/forx_xend200x_xloopexit_forx_xend200
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1074_if_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1074_if_link/if_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_34/forx_xbody193_forx_xend200x_xloopexit
      -- CP-element group 230: 	 branch_block_stmt_34/forx_xbody193_forx_xend200x_xloopexit_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_34/forx_xbody193_forx_xend200x_xloopexit_PhiReq/$exit
      -- CP-element group 230: 	 branch_block_stmt_34/merge_stmt_1080_PhiReqMerge
      -- CP-element group 230: 	 branch_block_stmt_34/merge_stmt_1080_PhiAck/$entry
      -- CP-element group 230: 	 branch_block_stmt_34/merge_stmt_1080_PhiAck/$exit
      -- CP-element group 230: 	 branch_block_stmt_34/merge_stmt_1080_PhiAck/dummy
      -- CP-element group 230: 	 branch_block_stmt_34/forx_xend200x_xloopexit_forx_xend200_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_34/forx_xend200x_xloopexit_forx_xend200_PhiReq/$exit
      -- 
    if_choice_transition_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1074_branch_ack_1, ack => testConfigure_CP_0_elements(230)); -- 
    -- CP-element group 231:  fork  transition  place  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	305 
    -- CP-element group 231: 	306 
    -- CP-element group 231:  members (12) 
      -- CP-element group 231: 	 branch_block_stmt_34/if_stmt_1074_else_link/$exit
      -- CP-element group 231: 	 branch_block_stmt_34/if_stmt_1074_else_link/else_choice_transition
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Sample/rr
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1074_branch_ack_0, ack => testConfigure_CP_0_elements(231)); -- 
    rr_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => type_cast_1049_inst_req_0); -- 
    cr_3227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => type_cast_1049_inst_req_1); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	310 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_Sample/ra
      -- 
    ra_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_0, ack => testConfigure_CP_0_elements(232)); -- 
    -- CP-element group 233:  transition  place  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	310 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (16) 
      -- CP-element group 233: 	 $exit
      -- CP-element group 233: 	 branch_block_stmt_34/$exit
      -- CP-element group 233: 	 branch_block_stmt_34/branch_block_stmt_34__exit__
      -- CP-element group 233: 	 branch_block_stmt_34/assign_stmt_1086__exit__
      -- CP-element group 233: 	 branch_block_stmt_34/return__
      -- CP-element group 233: 	 branch_block_stmt_34/merge_stmt_1088__exit__
      -- CP-element group 233: 	 branch_block_stmt_34/assign_stmt_1086/$exit
      -- CP-element group 233: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_Update/ca
      -- CP-element group 233: 	 branch_block_stmt_34/return___PhiReq/$entry
      -- CP-element group 233: 	 branch_block_stmt_34/return___PhiReq/$exit
      -- CP-element group 233: 	 branch_block_stmt_34/merge_stmt_1088_PhiReqMerge
      -- CP-element group 233: 	 branch_block_stmt_34/merge_stmt_1088_PhiAck/$entry
      -- CP-element group 233: 	 branch_block_stmt_34/merge_stmt_1088_PhiAck/$exit
      -- CP-element group 233: 	 branch_block_stmt_34/merge_stmt_1088_PhiAck/dummy
      -- 
    ca_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_1, ack => testConfigure_CP_0_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	32 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/Sample/ra
      -- 
    ra_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_78_inst_ack_0, ack => testConfigure_CP_0_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	32 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/Update/ca
      -- 
    ca_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_78_inst_ack_1, ack => testConfigure_CP_0_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	240 
    -- CP-element group 236:  members (5) 
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_78/SplitProtocol/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_req
      -- 
    phi_stmt_75_req_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_75_req_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(236), ack => phi_stmt_75_req_0); -- 
    testConfigure_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(234) & testConfigure_CP_0_elements(235);
      gj_testConfigure_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	32 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/Sample/ra
      -- 
    ra_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_0, ack => testConfigure_CP_0_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	32 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (2) 
      -- CP-element group 238: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/Update/ca
      -- 
    ca_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_1, ack => testConfigure_CP_0_elements(238)); -- 
    -- CP-element group 239:  join  transition  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (5) 
      -- CP-element group 239: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/$exit
      -- CP-element group 239: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/$exit
      -- CP-element group 239: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/$exit
      -- CP-element group 239: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_85/SplitProtocol/$exit
      -- CP-element group 239: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_req
      -- 
    phi_stmt_82_req_2693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_82_req_2693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(239), ack => phi_stmt_82_req_0); -- 
    testConfigure_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(237) & testConfigure_CP_0_elements(238);
      gj_testConfigure_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  join  transition  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	236 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	246 
    -- CP-element group 240:  members (1) 
      -- CP-element group 240: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(236) & testConfigure_CP_0_elements(239);
      gj_testConfigure_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  transition  output  delay-element  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	14 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	245 
    -- CP-element group 241:  members (4) 
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_75/$exit
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_sources/type_cast_81_konst_delay_trans
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_75/phi_stmt_75_req
      -- 
    phi_stmt_75_req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_75_req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => phi_stmt_75_req_1); -- 
    -- Element group testConfigure_CP_0_elements(241) is a control-delay.
    cp_element_241_delay: control_delay_element  generic map(name => " 241_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(14), ack => testConfigure_CP_0_elements(241), clk => clk, reset =>reset);
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	14 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/Sample/ra
      -- 
    ra_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_87_inst_ack_0, ack => testConfigure_CP_0_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	14 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/Update/ca
      -- 
    ca_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_87_inst_ack_1, ack => testConfigure_CP_0_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (5) 
      -- CP-element group 244: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/$exit
      -- CP-element group 244: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/$exit
      -- CP-element group 244: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/$exit
      -- CP-element group 244: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_sources/type_cast_87/SplitProtocol/$exit
      -- CP-element group 244: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_82/phi_stmt_82_req
      -- 
    phi_stmt_82_req_2727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_82_req_2727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => phi_stmt_82_req_1); -- 
    testConfigure_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(242) & testConfigure_CP_0_elements(243);
      gj_testConfigure_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	241 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (1) 
      -- CP-element group 245: 	 branch_block_stmt_34/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(241) & testConfigure_CP_0_elements(244);
      gj_testConfigure_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  merge  fork  transition  place  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	240 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_34/merge_stmt_74_PhiReqMerge
      -- CP-element group 246: 	 branch_block_stmt_34/merge_stmt_74_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(246) <= OrReduce(testConfigure_CP_0_elements(240) & testConfigure_CP_0_elements(245));
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (1) 
      -- CP-element group 247: 	 branch_block_stmt_34/merge_stmt_74_PhiAck/phi_stmt_75_ack
      -- 
    phi_stmt_75_ack_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_75_ack_0, ack => testConfigure_CP_0_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (1) 
      -- CP-element group 248: 	 branch_block_stmt_34/merge_stmt_74_PhiAck/phi_stmt_82_ack
      -- 
    phi_stmt_82_ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_82_ack_0, ack => testConfigure_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  fork  transition  place  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	26 
    -- CP-element group 249: 	29 
    -- CP-element group 249: 	15 
    -- CP-element group 249: 	16 
    -- CP-element group 249: 	17 
    -- CP-element group 249: 	18 
    -- CP-element group 249: 	20 
    -- CP-element group 249: 	22 
    -- CP-element group 249: 	23 
    -- CP-element group 249: 	25 
    -- CP-element group 249:  members (61) 
      -- CP-element group 249: 	 branch_block_stmt_34/merge_stmt_74__exit__
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137__entry__
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_update_start_
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_word_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_root_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_address_resized
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_update_start_
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_97_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_update_start_
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_resized_1
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_scaled_1
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_computed_1
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_resize_1/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_resize_1/$exit
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_resize_1/index_resize_req
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_resize_1/index_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_scale_1/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_scale_1/$exit
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_scale_1/scale_rename_req
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_index_scale_1/scale_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_update_start
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_Sample/req
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/array_obj_ref_103_final_index_sum_regn_Update/req
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/addr_of_104_complete/req
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_update_start_
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Update/word_access_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Update/word_access_complete/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_107_Update/word_access_complete/word_0/cr
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_addr_resize/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_addr_resize/$exit
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_addr_resize/base_resize_req
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_addr_resize/base_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_plus_offset/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_plus_offset/$exit
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_plus_offset/sum_rename_req
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_base_plus_offset/sum_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_word_addrgen/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_word_addrgen/$exit
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_word_addrgen/root_register_req
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_word_addrgen/root_register_ack
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/word_access_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/word_access_complete/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/ptr_deref_124_Update/word_access_complete/word_0/cr
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/RPIPE_ConvTranspose_input_pipe_132_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_update_start_
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_34/assign_stmt_94_to_assign_stmt_137/type_cast_136_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_34/merge_stmt_74_PhiAck/$exit
      -- 
    rr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_97_inst_req_0); -- 
    cr_251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_97_inst_req_1); -- 
    req_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => array_obj_ref_103_index_offset_req_0); -- 
    req_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => array_obj_ref_103_index_offset_req_1); -- 
    req_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => addr_of_104_final_reg_req_1); -- 
    cr_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => ptr_deref_107_store_0_req_1); -- 
    cr_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => ptr_deref_124_load_0_req_1); -- 
    rr_406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => RPIPE_ConvTranspose_input_pipe_132_inst_req_0); -- 
    cr_425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_136_inst_req_1); -- 
    testConfigure_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(247) & testConfigure_CP_0_elements(248);
      gj_testConfigure_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	33 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/Sample/ra
      -- 
    ra_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_148_inst_ack_0, ack => testConfigure_CP_0_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	33 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/Update/ca
      -- 
    ca_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_148_inst_ack_1, ack => testConfigure_CP_0_elements(251)); -- 
    -- CP-element group 252:  join  transition  place  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (8) 
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_sources/type_cast_148/SplitProtocol/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_145/phi_stmt_145_req
      -- CP-element group 252: 	 branch_block_stmt_34/merge_stmt_144_PhiReqMerge
      -- CP-element group 252: 	 branch_block_stmt_34/merge_stmt_144_PhiAck/$entry
      -- 
    phi_stmt_145_req_2763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_145_req_2763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(252), ack => phi_stmt_145_req_0); -- 
    testConfigure_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(250) & testConfigure_CP_0_elements(251);
      gj_testConfigure_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	257 
    -- CP-element group 253: 	258 
    -- CP-element group 253:  members (13) 
      -- CP-element group 253: 	 branch_block_stmt_34/merge_stmt_144__exit__
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend
      -- CP-element group 253: 	 branch_block_stmt_34/merge_stmt_144_PhiAck/$exit
      -- CP-element group 253: 	 branch_block_stmt_34/merge_stmt_144_PhiAck/phi_stmt_145_ack
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/Sample/rr
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/Update/cr
      -- 
    phi_stmt_145_ack_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_145_ack_0, ack => testConfigure_CP_0_elements(253)); -- 
    rr_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => type_cast_157_inst_req_0); -- 
    cr_2818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => type_cast_157_inst_req_1); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	13 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/Sample/ra
      -- 
    ra_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_0, ack => testConfigure_CP_0_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	13 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (2) 
      -- CP-element group 255: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/Update/ca
      -- 
    ca_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_1, ack => testConfigure_CP_0_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	260 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/$exit
      -- CP-element group 256: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/$exit
      -- CP-element group 256: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/$exit
      -- CP-element group 256: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/$exit
      -- CP-element group 256: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_155/SplitProtocol/$exit
      -- CP-element group 256: 	 branch_block_stmt_34/entry_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_req
      -- 
    phi_stmt_152_req_2794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_152_req_2794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(256), ack => phi_stmt_152_req_0); -- 
    testConfigure_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(254) & testConfigure_CP_0_elements(255);
      gj_testConfigure_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	253 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (2) 
      -- CP-element group 257: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/Sample/ra
      -- 
    ra_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_0, ack => testConfigure_CP_0_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	253 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/Update/ca
      -- 
    ca_2819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_1, ack => testConfigure_CP_0_elements(258)); -- 
    -- CP-element group 259:  join  transition  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 259: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/$exit
      -- CP-element group 259: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/$exit
      -- CP-element group 259: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/$exit
      -- CP-element group 259: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_sources/type_cast_157/SplitProtocol/$exit
      -- CP-element group 259: 	 branch_block_stmt_34/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_152/phi_stmt_152_req
      -- 
    phi_stmt_152_req_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_152_req_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => phi_stmt_152_req_1); -- 
    testConfigure_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(257) & testConfigure_CP_0_elements(258);
      gj_testConfigure_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  merge  transition  place  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	256 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (2) 
      -- CP-element group 260: 	 branch_block_stmt_34/merge_stmt_151_PhiReqMerge
      -- CP-element group 260: 	 branch_block_stmt_34/merge_stmt_151_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(260) <= OrReduce(testConfigure_CP_0_elements(256) & testConfigure_CP_0_elements(259));
    -- CP-element group 261:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	34 
    -- CP-element group 261: 	35 
    -- CP-element group 261:  members (35) 
      -- CP-element group 261: 	 branch_block_stmt_34/merge_stmt_151__exit__
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174__entry__
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_update_start_
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_word_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_root_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_address_resized
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_addr_resize/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_addr_resize/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_addr_resize/base_resize_req
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_addr_resize/base_resize_ack
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_plus_offset/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_plus_offset/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_plus_offset/sum_rename_req
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_base_plus_offset/sum_rename_ack
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_word_addrgen/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_word_addrgen/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_word_addrgen/root_register_req
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_word_addrgen/root_register_ack
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/ptr_deref_166_Split/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/ptr_deref_166_Split/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/ptr_deref_166_Split/split_req
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/ptr_deref_166_Split/split_ack
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/word_access_start/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/word_access_start/word_0/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Sample/word_access_start/word_0/rr
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Update/word_access_complete/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Update/word_access_complete/word_0/$entry
      -- CP-element group 261: 	 branch_block_stmt_34/assign_stmt_164_to_assign_stmt_174/ptr_deref_166_Update/word_access_complete/word_0/cr
      -- CP-element group 261: 	 branch_block_stmt_34/merge_stmt_151_PhiAck/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/merge_stmt_151_PhiAck/phi_stmt_152_ack
      -- 
    phi_stmt_152_ack_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_152_ack_0, ack => testConfigure_CP_0_elements(261)); -- 
    rr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(261), ack => ptr_deref_166_store_0_req_0); -- 
    cr_498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(261), ack => ptr_deref_166_store_0_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	56 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (2) 
      -- CP-element group 262: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/Sample/ra
      -- 
    ra_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_187_inst_ack_0, ack => testConfigure_CP_0_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	56 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (2) 
      -- CP-element group 263: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/Update/ca
      -- 
    ca_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_187_inst_ack_1, ack => testConfigure_CP_0_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/$exit
      -- CP-element group 264: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/$exit
      -- CP-element group 264: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/$exit
      -- CP-element group 264: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/$exit
      -- CP-element group 264: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_187/SplitProtocol/$exit
      -- CP-element group 264: 	 branch_block_stmt_34/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_req
      -- 
    phi_stmt_184_req_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_184_req_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => phi_stmt_184_req_0); -- 
    testConfigure_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(262) & testConfigure_CP_0_elements(263);
      gj_testConfigure_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  transition  output  delay-element  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	37 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (5) 
      -- CP-element group 265: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/$exit
      -- CP-element group 265: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_184/$exit
      -- CP-element group 265: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/$exit
      -- CP-element group 265: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_sources/type_cast_190_konst_delay_trans
      -- CP-element group 265: 	 branch_block_stmt_34/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_184/phi_stmt_184_req
      -- 
    phi_stmt_184_req_2874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_184_req_2874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(265), ack => phi_stmt_184_req_1); -- 
    -- Element group testConfigure_CP_0_elements(265) is a control-delay.
    cp_element_265_delay: control_delay_element  generic map(name => " 265_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(37), ack => testConfigure_CP_0_elements(265), clk => clk, reset =>reset);
    -- CP-element group 266:  merge  transition  place  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_34/merge_stmt_183_PhiReqMerge
      -- CP-element group 266: 	 branch_block_stmt_34/merge_stmt_183_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(266) <= OrReduce(testConfigure_CP_0_elements(264) & testConfigure_CP_0_elements(265));
    -- CP-element group 267:  fork  transition  place  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	38 
    -- CP-element group 267: 	39 
    -- CP-element group 267: 	40 
    -- CP-element group 267: 	41 
    -- CP-element group 267: 	43 
    -- CP-element group 267: 	44 
    -- CP-element group 267: 	47 
    -- CP-element group 267: 	50 
    -- CP-element group 267: 	51 
    -- CP-element group 267: 	53 
    -- CP-element group 267:  members (62) 
      -- CP-element group 267: 	 branch_block_stmt_34/merge_stmt_183__exit__
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240__entry__
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_update_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_200_Update/cr
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_update_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_resized_1
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_scaled_1
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_computed_1
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_resize_1/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_resize_1/$exit
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_resize_1/index_resize_req
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_resize_1/index_resize_ack
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_scale_1/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_scale_1/$exit
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_scale_1/scale_rename_req
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_index_scale_1/scale_rename_ack
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_update_start
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_Sample/req
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/array_obj_ref_206_final_index_sum_regn_Update/req
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/addr_of_207_complete/req
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/RPIPE_ConvTranspose_input_pipe_210_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_update_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/type_cast_214_Update/cr
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_update_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Update/word_access_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Update/word_access_complete/word_0/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_217_Update/word_access_complete/word_0/cr
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_update_start_
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_word_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_root_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_address_resized
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_addr_resize/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_addr_resize/$exit
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_addr_resize/base_resize_req
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_addr_resize/base_resize_ack
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_plus_offset/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_plus_offset/$exit
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_plus_offset/sum_rename_req
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_base_plus_offset/sum_rename_ack
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_word_addrgen/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_word_addrgen/$exit
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_word_addrgen/root_register_req
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_word_addrgen/root_register_ack
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/word_access_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/word_access_complete/word_0/$entry
      -- CP-element group 267: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_240/ptr_deref_234_Update/word_access_complete/word_0/cr
      -- CP-element group 267: 	 branch_block_stmt_34/merge_stmt_183_PhiAck/$exit
      -- CP-element group 267: 	 branch_block_stmt_34/merge_stmt_183_PhiAck/phi_stmt_184_ack
      -- 
    phi_stmt_184_ack_2879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_184_ack_0, ack => testConfigure_CP_0_elements(267)); -- 
    rr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_200_inst_req_0); -- 
    cr_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_200_inst_req_1); -- 
    req_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => array_obj_ref_206_index_offset_req_0); -- 
    req_565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => array_obj_ref_206_index_offset_req_1); -- 
    req_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => addr_of_207_final_reg_req_1); -- 
    rr_589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => RPIPE_ConvTranspose_input_pipe_210_inst_req_0); -- 
    cr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_214_inst_req_1); -- 
    cr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => ptr_deref_217_store_0_req_1); -- 
    cr_703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => ptr_deref_234_load_0_req_1); -- 
    -- CP-element group 268:  merge  fork  transition  place  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	36 
    -- CP-element group 268: 	57 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	58 
    -- CP-element group 268: 	61 
    -- CP-element group 268:  members (13) 
      -- CP-element group 268: 	 branch_block_stmt_34/merge_stmt_249__exit__
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256__entry__
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/$entry
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/RPIPE_ConvTranspose_input_pipe_251_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_update_start_
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_34/assign_stmt_252_to_assign_stmt_256/type_cast_255_Update/cr
      -- CP-element group 268: 	 branch_block_stmt_34/merge_stmt_249_PhiReqMerge
      -- CP-element group 268: 	 branch_block_stmt_34/merge_stmt_249_PhiAck/$entry
      -- CP-element group 268: 	 branch_block_stmt_34/merge_stmt_249_PhiAck/$exit
      -- CP-element group 268: 	 branch_block_stmt_34/merge_stmt_249_PhiAck/dummy
      -- 
    rr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(268), ack => RPIPE_ConvTranspose_input_pipe_251_inst_req_0); -- 
    cr_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(268), ack => type_cast_255_inst_req_1); -- 
    testConfigure_CP_0_elements(268) <= OrReduce(testConfigure_CP_0_elements(36) & testConfigure_CP_0_elements(57));
    -- CP-element group 269:  transition  output  delay-element  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	61 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	273 
    -- CP-element group 269:  members (4) 
      -- CP-element group 269: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_259/$exit
      -- CP-element group 269: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/$exit
      -- CP-element group 269: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_263_konst_delay_trans
      -- CP-element group 269: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_req
      -- 
    phi_stmt_259_req_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_259_req_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(269), ack => phi_stmt_259_req_0); -- 
    -- Element group testConfigure_CP_0_elements(269) is a control-delay.
    cp_element_269_delay: control_delay_element  generic map(name => " 269_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(61), ack => testConfigure_CP_0_elements(269), clk => clk, reset =>reset);
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	61 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/Sample/ra
      -- 
    ra_2930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_0, ack => testConfigure_CP_0_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	61 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (2) 
      -- CP-element group 271: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/Update/ca
      -- 
    ca_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_1, ack => testConfigure_CP_0_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (5) 
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/$exit
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/$exit
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/$exit
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_269/SplitProtocol/$exit
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_req
      -- 
    phi_stmt_266_req_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_266_req_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => phi_stmt_266_req_0); -- 
    testConfigure_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(270) & testConfigure_CP_0_elements(271);
      gj_testConfigure_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	269 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	281 
    -- CP-element group 273:  members (1) 
      -- CP-element group 273: 	 branch_block_stmt_34/bbx_xnph221_forx_xbody28_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(269) & testConfigure_CP_0_elements(272);
      gj_testConfigure_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	72 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/Sample/ra
      -- 
    ra_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_0, ack => testConfigure_CP_0_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	72 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (2) 
      -- CP-element group 275: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/Update/ca
      -- 
    ca_2961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_1, ack => testConfigure_CP_0_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	280 
    -- CP-element group 276:  members (5) 
      -- CP-element group 276: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/$exit
      -- CP-element group 276: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/$exit
      -- CP-element group 276: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/$exit
      -- CP-element group 276: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_sources/type_cast_265/SplitProtocol/$exit
      -- CP-element group 276: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_259/phi_stmt_259_req
      -- 
    phi_stmt_259_req_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_259_req_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => phi_stmt_259_req_1); -- 
    testConfigure_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(274) & testConfigure_CP_0_elements(275);
      gj_testConfigure_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	72 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (2) 
      -- CP-element group 277: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/Sample/ra
      -- 
    ra_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_271_inst_ack_0, ack => testConfigure_CP_0_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	72 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/Update/ca
      -- 
    ca_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_271_inst_ack_1, ack => testConfigure_CP_0_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (5) 
      -- CP-element group 279: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_sources/type_cast_271/SplitProtocol/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_266/phi_stmt_266_req
      -- 
    phi_stmt_266_req_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_266_req_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => phi_stmt_266_req_1); -- 
    testConfigure_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(277) & testConfigure_CP_0_elements(278);
      gj_testConfigure_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  join  transition  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	276 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_34/forx_xbody28_forx_xbody28_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(276) & testConfigure_CP_0_elements(279);
      gj_testConfigure_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  merge  fork  transition  place  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	273 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_34/merge_stmt_258_PhiReqMerge
      -- CP-element group 281: 	 branch_block_stmt_34/merge_stmt_258_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(281) <= OrReduce(testConfigure_CP_0_elements(273) & testConfigure_CP_0_elements(280));
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_34/merge_stmt_258_PhiAck/phi_stmt_259_ack
      -- 
    phi_stmt_259_ack_2990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_259_ack_0, ack => testConfigure_CP_0_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_34/merge_stmt_258_PhiAck/phi_stmt_266_ack
      -- 
    phi_stmt_266_ack_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_266_ack_0, ack => testConfigure_CP_0_elements(283)); -- 
    -- CP-element group 284:  join  fork  transition  place  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	62 
    -- CP-element group 284: 	63 
    -- CP-element group 284: 	65 
    -- CP-element group 284: 	66 
    -- CP-element group 284: 	69 
    -- CP-element group 284:  members (42) 
      -- CP-element group 284: 	 branch_block_stmt_34/merge_stmt_258__exit__
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300__entry__
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_final_index_sum_regn/ack
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_request/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_request/req
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_complete/req
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_update_start_
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/addr_of_276_update_start_
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_offset_calculated
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_resized_0
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_scaled_0
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_computed_0
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_resize_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_resize_0/$exit
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_resize_0/index_resize_req
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_resize_0/index_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_scale_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_scale_0/$exit
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_scale_0/scale_rename_req
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_index_scale_0/scale_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_final_index_sum_regn/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_final_index_sum_regn/$exit
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/array_obj_ref_275_final_index_sum_regn/req
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/ptr_deref_279_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/RPIPE_ConvTranspose_input_pipe_283_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_update_start_
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_34/assign_stmt_277_to_assign_stmt_300/type_cast_287_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_34/merge_stmt_258_PhiAck/$exit
      -- 
    req_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => addr_of_276_final_reg_req_0); -- 
    req_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => addr_of_276_final_reg_req_1); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => ptr_deref_279_store_0_req_1); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => RPIPE_ConvTranspose_input_pipe_283_inst_req_0); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => type_cast_287_inst_req_1); -- 
    testConfigure_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(282) & testConfigure_CP_0_elements(283);
      gj_testConfigure_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	71 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/Sample/ra
      -- 
    ra_3015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_0, ack => testConfigure_CP_0_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	71 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/Update/ca
      -- 
    ca_3020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_1, ack => testConfigure_CP_0_elements(286)); -- 
    -- CP-element group 287:  join  transition  place  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (8) 
      -- CP-element group 287: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/$exit
      -- CP-element group 287: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/$exit
      -- CP-element group 287: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/$exit
      -- CP-element group 287: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/$exit
      -- CP-element group 287: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_sources/type_cast_311/SplitProtocol/$exit
      -- CP-element group 287: 	 branch_block_stmt_34/forx_xbody28_forx_xend37_PhiReq/phi_stmt_308/phi_stmt_308_req
      -- CP-element group 287: 	 branch_block_stmt_34/merge_stmt_307_PhiReqMerge
      -- CP-element group 287: 	 branch_block_stmt_34/merge_stmt_307_PhiAck/$entry
      -- 
    phi_stmt_308_req_3021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_308_req_3021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => phi_stmt_308_req_0); -- 
    testConfigure_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(285) & testConfigure_CP_0_elements(286);
      gj_testConfigure_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  merge  transition  place  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	73 
    -- CP-element group 288:  members (4) 
      -- CP-element group 288: 	 branch_block_stmt_34/merge_stmt_307__exit__
      -- CP-element group 288: 	 branch_block_stmt_34/assign_stmt_315_to_assign_stmt_501__entry__
      -- CP-element group 288: 	 branch_block_stmt_34/merge_stmt_307_PhiAck/$exit
      -- CP-element group 288: 	 branch_block_stmt_34/merge_stmt_307_PhiAck/phi_stmt_308_ack
      -- 
    phi_stmt_308_ack_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_308_ack_0, ack => testConfigure_CP_0_elements(288)); -- 
    -- CP-element group 289:  merge  branch  transition  place  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	120 
    -- CP-element group 289: 	166 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	122 
    -- CP-element group 289: 	123 
    -- CP-element group 289:  members (17) 
      -- CP-element group 289: 	 branch_block_stmt_34/merge_stmt_510__exit__
      -- CP-element group 289: 	 branch_block_stmt_34/assign_stmt_516_to_assign_stmt_522__entry__
      -- CP-element group 289: 	 branch_block_stmt_34/assign_stmt_516_to_assign_stmt_522__exit__
      -- CP-element group 289: 	 branch_block_stmt_34/if_stmt_523__entry__
      -- CP-element group 289: 	 branch_block_stmt_34/assign_stmt_516_to_assign_stmt_522/$entry
      -- CP-element group 289: 	 branch_block_stmt_34/assign_stmt_516_to_assign_stmt_522/$exit
      -- CP-element group 289: 	 branch_block_stmt_34/if_stmt_523_dead_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_34/if_stmt_523_eval_test/$entry
      -- CP-element group 289: 	 branch_block_stmt_34/if_stmt_523_eval_test/$exit
      -- CP-element group 289: 	 branch_block_stmt_34/if_stmt_523_eval_test/branch_req
      -- CP-element group 289: 	 branch_block_stmt_34/R_cmp124208_524_place
      -- CP-element group 289: 	 branch_block_stmt_34/if_stmt_523_if_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_34/if_stmt_523_else_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_34/merge_stmt_510_PhiReqMerge
      -- CP-element group 289: 	 branch_block_stmt_34/merge_stmt_510_PhiAck/$entry
      -- CP-element group 289: 	 branch_block_stmt_34/merge_stmt_510_PhiAck/$exit
      -- CP-element group 289: 	 branch_block_stmt_34/merge_stmt_510_PhiAck/dummy
      -- 
    branch_req_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => if_stmt_523_branch_req_0); -- 
    testConfigure_CP_0_elements(289) <= OrReduce(testConfigure_CP_0_elements(120) & testConfigure_CP_0_elements(166));
    -- CP-element group 290:  transition  output  delay-element  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	125 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	294 
    -- CP-element group 290:  members (5) 
      -- CP-element group 290: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67_PhiReq/$exit
      -- CP-element group 290: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_565/$exit
      -- CP-element group 290: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/$exit
      -- CP-element group 290: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_569_konst_delay_trans
      -- CP-element group 290: 	 branch_block_stmt_34/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_req
      -- 
    phi_stmt_565_req_3072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_565_req_3072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(290), ack => phi_stmt_565_req_0); -- 
    -- Element group testConfigure_CP_0_elements(290) is a control-delay.
    cp_element_290_delay: control_delay_element  generic map(name => " 290_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(125), ack => testConfigure_CP_0_elements(290), clk => clk, reset =>reset);
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	167 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (2) 
      -- CP-element group 291: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/Sample/ra
      -- 
    ra_3092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_571_inst_ack_0, ack => testConfigure_CP_0_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	167 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (2) 
      -- CP-element group 292: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/Update/ca
      -- 
    ca_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_571_inst_ack_1, ack => testConfigure_CP_0_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/$exit
      -- CP-element group 293: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/$exit
      -- CP-element group 293: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/$exit
      -- CP-element group 293: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/$exit
      -- CP-element group 293: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_sources/type_cast_571/SplitProtocol/$exit
      -- CP-element group 293: 	 branch_block_stmt_34/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_565/phi_stmt_565_req
      -- 
    phi_stmt_565_req_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_565_req_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => phi_stmt_565_req_1); -- 
    testConfigure_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(291) & testConfigure_CP_0_elements(292);
      gj_testConfigure_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  merge  transition  place  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	290 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (2) 
      -- CP-element group 294: 	 branch_block_stmt_34/merge_stmt_564_PhiReqMerge
      -- CP-element group 294: 	 branch_block_stmt_34/merge_stmt_564_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(294) <= OrReduce(testConfigure_CP_0_elements(290) & testConfigure_CP_0_elements(293));
    -- CP-element group 295:  fork  transition  place  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	126 
    -- CP-element group 295: 	127 
    -- CP-element group 295: 	129 
    -- CP-element group 295: 	130 
    -- CP-element group 295: 	133 
    -- CP-element group 295: 	137 
    -- CP-element group 295: 	141 
    -- CP-element group 295: 	145 
    -- CP-element group 295: 	149 
    -- CP-element group 295: 	153 
    -- CP-element group 295: 	157 
    -- CP-element group 295: 	161 
    -- CP-element group 295: 	164 
    -- CP-element group 295:  members (56) 
      -- CP-element group 295: 	 branch_block_stmt_34/merge_stmt_564__exit__
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727__entry__
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_resized_1
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_scaled_1
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_computed_1
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_resize_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_resize_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_resize_1/index_resize_req
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_resize_1/index_resize_ack
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_scale_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_scale_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_scale_1/scale_rename_req
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_index_scale_1/scale_rename_ack
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_update_start
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_Sample/req
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/array_obj_ref_577_final_index_sum_regn_Update/req
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/addr_of_578_complete/req
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/RPIPE_ConvTranspose_input_pipe_581_Sample/rr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_585_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_598_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_616_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_634_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_652_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_670_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_688_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/type_cast_706_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_update_start_
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Update/word_access_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Update/word_access_complete/word_0/$entry
      -- CP-element group 295: 	 branch_block_stmt_34/assign_stmt_579_to_assign_stmt_727/ptr_deref_714_Update/word_access_complete/word_0/cr
      -- CP-element group 295: 	 branch_block_stmt_34/merge_stmt_564_PhiAck/$exit
      -- CP-element group 295: 	 branch_block_stmt_34/merge_stmt_564_PhiAck/phi_stmt_565_ack
      -- 
    phi_stmt_565_ack_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_565_ack_0, ack => testConfigure_CP_0_elements(295)); -- 
    req_1635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => array_obj_ref_577_index_offset_req_0); -- 
    req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => array_obj_ref_577_index_offset_req_1); -- 
    req_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => addr_of_578_final_reg_req_1); -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => RPIPE_ConvTranspose_input_pipe_581_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_585_inst_req_1); -- 
    cr_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_598_inst_req_1); -- 
    cr_1739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_616_inst_req_1); -- 
    cr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_634_inst_req_1); -- 
    cr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_652_inst_req_1); -- 
    cr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_670_inst_req_1); -- 
    cr_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_688_inst_req_1); -- 
    cr_1879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_706_inst_req_1); -- 
    cr_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => ptr_deref_714_store_0_req_1); -- 
    -- CP-element group 296:  transition  output  delay-element  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	169 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	300 
    -- CP-element group 296:  members (5) 
      -- CP-element group 296: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126_PhiReq/$exit
      -- CP-element group 296: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_775/$exit
      -- CP-element group 296: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/$exit
      -- CP-element group 296: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_779_konst_delay_trans
      -- CP-element group 296: 	 branch_block_stmt_34/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_req
      -- 
    phi_stmt_775_req_3126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_775_req_3126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(296), ack => phi_stmt_775_req_0); -- 
    -- Element group testConfigure_CP_0_elements(296) is a control-delay.
    cp_element_296_delay: control_delay_element  generic map(name => " 296_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(169), ack => testConfigure_CP_0_elements(296), clk => clk, reset =>reset);
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	211 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (2) 
      -- CP-element group 297: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/Sample/ra
      -- 
    ra_3146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_0, ack => testConfigure_CP_0_elements(297)); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	211 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (2) 
      -- CP-element group 298: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/Update/ca
      -- 
    ca_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_1, ack => testConfigure_CP_0_elements(298)); -- 
    -- CP-element group 299:  join  transition  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/$exit
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/$exit
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/$exit
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/$exit
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_sources/type_cast_781/SplitProtocol/$exit
      -- CP-element group 299: 	 branch_block_stmt_34/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_775/phi_stmt_775_req
      -- 
    phi_stmt_775_req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_775_req_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(299), ack => phi_stmt_775_req_1); -- 
    testConfigure_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(297) & testConfigure_CP_0_elements(298);
      gj_testConfigure_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  merge  transition  place  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	296 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (2) 
      -- CP-element group 300: 	 branch_block_stmt_34/merge_stmt_774_PhiReqMerge
      -- CP-element group 300: 	 branch_block_stmt_34/merge_stmt_774_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(300) <= OrReduce(testConfigure_CP_0_elements(296) & testConfigure_CP_0_elements(299));
    -- CP-element group 301:  fork  transition  place  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	170 
    -- CP-element group 301: 	171 
    -- CP-element group 301: 	173 
    -- CP-element group 301: 	174 
    -- CP-element group 301: 	177 
    -- CP-element group 301: 	181 
    -- CP-element group 301: 	185 
    -- CP-element group 301: 	189 
    -- CP-element group 301: 	193 
    -- CP-element group 301: 	197 
    -- CP-element group 301: 	201 
    -- CP-element group 301: 	205 
    -- CP-element group 301: 	208 
    -- CP-element group 301:  members (56) 
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_34/merge_stmt_774__exit__
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937__entry__
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_862_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_898_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Update/word_access_complete/word_0/cr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Update/word_access_complete/word_0/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Update/word_access_complete/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/ptr_deref_924_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_916_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_880_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_resized_1
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_scaled_1
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_computed_1
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_resize_1/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_resize_1/$exit
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_resize_1/index_resize_req
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_resize_1/index_resize_ack
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_scale_1/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_scale_1/$exit
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_scale_1/scale_rename_req
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_index_scale_1/scale_rename_ack
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_update_start
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_Sample/req
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/array_obj_ref_787_final_index_sum_regn_Update/req
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_complete/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/addr_of_788_complete/req
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/RPIPE_ConvTranspose_input_pipe_791_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_795_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_808_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_826_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_34/assign_stmt_789_to_assign_stmt_937/type_cast_844_update_start_
      -- CP-element group 301: 	 branch_block_stmt_34/merge_stmt_774_PhiAck/$exit
      -- CP-element group 301: 	 branch_block_stmt_34/merge_stmt_774_PhiAck/phi_stmt_775_ack
      -- 
    phi_stmt_775_ack_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_775_ack_0, ack => testConfigure_CP_0_elements(301)); -- 
    cr_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_898_inst_req_1); -- 
    cr_2154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_862_inst_req_1); -- 
    cr_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_916_inst_req_1); -- 
    cr_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => ptr_deref_924_store_0_req_1); -- 
    cr_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_844_inst_req_1); -- 
    cr_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_880_inst_req_1); -- 
    req_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => array_obj_ref_787_index_offset_req_0); -- 
    req_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => array_obj_ref_787_index_offset_req_1); -- 
    req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => addr_of_788_final_reg_req_1); -- 
    rr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => RPIPE_ConvTranspose_input_pipe_791_inst_req_0); -- 
    cr_2042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_795_inst_req_1); -- 
    cr_2070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_808_inst_req_1); -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_826_inst_req_1); -- 
    -- CP-element group 302:  merge  place  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	122 
    -- CP-element group 302: 	210 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (1) 
      -- CP-element group 302: 	 branch_block_stmt_34/merge_stmt_946_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(302) <= OrReduce(testConfigure_CP_0_elements(122) & testConfigure_CP_0_elements(210));
    -- CP-element group 303:  join  fork  transition  place  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	212 
    -- CP-element group 303: 	213 
    -- CP-element group 303: 	214 
    -- CP-element group 303: 	215 
    -- CP-element group 303: 	216 
    -- CP-element group 303: 	217 
    -- CP-element group 303:  members (84) 
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/merge_stmt_946__exit__
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998__entry__
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_update_start_
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_957_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_update_start_
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_981_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_update_start_
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_34/assign_stmt_954_to_assign_stmt_998/ptr_deref_969_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/merge_stmt_946_PhiAck/$entry
      -- CP-element group 303: 	 branch_block_stmt_34/merge_stmt_946_PhiAck/$exit
      -- CP-element group 303: 	 branch_block_stmt_34/merge_stmt_946_PhiAck/dummy
      -- 
    rr_2444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_981_load_0_req_0); -- 
    cr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_981_load_0_req_1); -- 
    rr_2344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_957_load_0_req_0); -- 
    cr_2355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_957_load_0_req_1); -- 
    rr_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_969_load_0_req_0); -- 
    cr_2405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_969_load_0_req_1); -- 
    testConfigure_CP_0_elements(303) <= testConfigure_CP_0_elements(302);
    -- CP-element group 304:  transition  output  delay-element  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	222 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	308 
    -- CP-element group 304:  members (5) 
      -- CP-element group 304: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193_PhiReq/$exit
      -- CP-element group 304: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1043/$exit
      -- CP-element group 304: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/$exit
      -- CP-element group 304: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1047_konst_delay_trans
      -- CP-element group 304: 	 branch_block_stmt_34/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_req
      -- 
    phi_stmt_1043_req_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1043_req_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(304), ack => phi_stmt_1043_req_0); -- 
    -- Element group testConfigure_CP_0_elements(304) is a control-delay.
    cp_element_304_delay: control_delay_element  generic map(name => " 304_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(222), ack => testConfigure_CP_0_elements(304), clk => clk, reset =>reset);
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	231 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Sample/ra
      -- 
    ra_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1049_inst_ack_0, ack => testConfigure_CP_0_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	231 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (2) 
      -- CP-element group 306: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/Update/ca
      -- 
    ca_3228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1049_inst_ack_1, ack => testConfigure_CP_0_elements(306)); -- 
    -- CP-element group 307:  join  transition  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/$exit
      -- CP-element group 307: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/$exit
      -- CP-element group 307: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/$exit
      -- CP-element group 307: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/$exit
      -- CP-element group 307: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_sources/type_cast_1049/SplitProtocol/$exit
      -- CP-element group 307: 	 branch_block_stmt_34/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1043/phi_stmt_1043_req
      -- 
    phi_stmt_1043_req_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1043_req_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(307), ack => phi_stmt_1043_req_1); -- 
    testConfigure_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(305) & testConfigure_CP_0_elements(306);
      gj_testConfigure_cp_element_group_307 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  merge  transition  place  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	304 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (2) 
      -- CP-element group 308: 	 branch_block_stmt_34/merge_stmt_1042_PhiReqMerge
      -- CP-element group 308: 	 branch_block_stmt_34/merge_stmt_1042_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(308) <= OrReduce(testConfigure_CP_0_elements(304) & testConfigure_CP_0_elements(307));
    -- CP-element group 309:  fork  transition  place  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	223 
    -- CP-element group 309: 	224 
    -- CP-element group 309: 	226 
    -- CP-element group 309: 	228 
    -- CP-element group 309:  members (29) 
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_resize_1/index_resize_ack
      -- CP-element group 309: 	 branch_block_stmt_34/merge_stmt_1042__exit__
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073__entry__
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_scale_1/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_scale_1/$exit
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_scale_1/scale_rename_req
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_scale_1/scale_rename_ack
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_resize_1/index_resize_req
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_resize_1/$exit
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_resize_1/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_computed_1
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_complete/req
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_Update/req
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_scaled_1
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_index_resized_1
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_complete/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_Sample/req
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/array_obj_ref_1055_final_index_sum_regn_update_start
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_update_start_
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/addr_of_1056_update_start_
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Update/word_access_complete/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Update/word_access_complete/word_0/$entry
      -- CP-element group 309: 	 branch_block_stmt_34/assign_stmt_1057_to_assign_stmt_1073/ptr_deref_1059_Update/word_access_complete/word_0/cr
      -- CP-element group 309: 	 branch_block_stmt_34/merge_stmt_1042_PhiAck/$exit
      -- CP-element group 309: 	 branch_block_stmt_34/merge_stmt_1042_PhiAck/phi_stmt_1043_ack
      -- 
    phi_stmt_1043_ack_3234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1043_ack_0, ack => testConfigure_CP_0_elements(309)); -- 
    req_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => addr_of_1056_final_reg_req_1); -- 
    req_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => array_obj_ref_1055_index_offset_req_1); -- 
    req_2525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => array_obj_ref_1055_index_offset_req_0); -- 
    cr_2595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => ptr_deref_1059_store_0_req_1); -- 
    -- CP-element group 310:  merge  fork  transition  place  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	220 
    -- CP-element group 310: 	230 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	232 
    -- CP-element group 310: 	233 
    -- CP-element group 310:  members (13) 
      -- CP-element group 310: 	 branch_block_stmt_34/merge_stmt_1082__exit__
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1086__entry__
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1086/$entry
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_update_start_
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_Sample/rr
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_34/assign_stmt_1086/type_cast_1085_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_34/merge_stmt_1082_PhiReqMerge
      -- CP-element group 310: 	 branch_block_stmt_34/merge_stmt_1082_PhiAck/$entry
      -- CP-element group 310: 	 branch_block_stmt_34/merge_stmt_1082_PhiAck/$exit
      -- CP-element group 310: 	 branch_block_stmt_34/merge_stmt_1082_PhiAck/dummy
      -- 
    rr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(310), ack => type_cast_1085_inst_req_0); -- 
    cr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(310), ack => type_cast_1085_inst_req_1); -- 
    testConfigure_CP_0_elements(310) <= OrReduce(testConfigure_CP_0_elements(220) & testConfigure_CP_0_elements(230));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar240_786_resized : std_logic_vector(10 downto 0);
    signal R_indvar240_786_scaled : std_logic_vector(10 downto 0);
    signal R_indvar250_576_resized : std_logic_vector(13 downto 0);
    signal R_indvar250_576_scaled : std_logic_vector(13 downto 0);
    signal R_indvar260_274_resized : std_logic_vector(0 downto 0);
    signal R_indvar260_274_scaled : std_logic_vector(0 downto 0);
    signal R_indvar263_205_resized : std_logic_vector(6 downto 0);
    signal R_indvar263_205_scaled : std_logic_vector(6 downto 0);
    signal R_indvar268_102_resized : std_logic_vector(6 downto 0);
    signal R_indvar268_102_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_1054_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1054_scaled : std_logic_vector(13 downto 0);
    signal STORE_padding_313_data_0 : std_logic_vector(15 downto 0);
    signal STORE_padding_313_word_address_0 : std_logic_vector(0 downto 0);
    signal add104_694 : std_logic_vector(63 downto 0);
    signal add110_712 : std_logic_vector(63 downto 0);
    signal add136_814 : std_logic_vector(63 downto 0);
    signal add142_832 : std_logic_vector(63 downto 0);
    signal add148_850 : std_logic_vector(63 downto 0);
    signal add154_868 : std_logic_vector(63 downto 0);
    signal add160_886 : std_logic_vector(63 downto 0);
    signal add166_904 : std_logic_vector(63 downto 0);
    signal add172_922 : std_logic_vector(63 downto 0);
    signal add80_622 : std_logic_vector(63 downto 0);
    signal add86_640 : std_logic_vector(63 downto 0);
    signal add92_658 : std_logic_vector(63 downto 0);
    signal add98_676 : std_logic_vector(63 downto 0);
    signal add_604 : std_logic_vector(63 downto 0);
    signal array_obj_ref_103_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_103_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_103_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_103_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_103_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_103_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1055_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1055_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_206_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_206_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_206_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_206_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_206_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_206_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_275_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_275_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_275_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_275_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_577_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_577_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_577_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_577_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_577_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_577_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_787_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_787_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_787_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_787_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_787_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_787_root_address : std_logic_vector(10 downto 0);
    signal arrayidx114_579 : std_logic_vector(31 downto 0);
    signal arrayidx176_789 : std_logic_vector(31 downto 0);
    signal arrayidx196_1057 : std_logic_vector(31 downto 0);
    signal arrayidx19_208 : std_logic_vector(31 downto 0);
    signal arrayidx33_277 : std_logic_vector(31 downto 0);
    signal arrayidx_105 : std_logic_vector(31 downto 0);
    signal call101_685 : std_logic_vector(7 downto 0);
    signal call107_703 : std_logic_vector(7 downto 0);
    signal call129_792 : std_logic_vector(7 downto 0);
    signal call133_805 : std_logic_vector(7 downto 0);
    signal call139_823 : std_logic_vector(7 downto 0);
    signal call145_841 : std_logic_vector(7 downto 0);
    signal call151_859 : std_logic_vector(7 downto 0);
    signal call157_877 : std_logic_vector(7 downto 0);
    signal call15_211 : std_logic_vector(7 downto 0);
    signal call163_895 : std_logic_vector(7 downto 0);
    signal call169_913 : std_logic_vector(7 downto 0);
    signal call29217_252 : std_logic_vector(7 downto 0);
    signal call29_284 : std_logic_vector(7 downto 0);
    signal call3228_61 : std_logic_vector(7 downto 0);
    signal call3_133 : std_logic_vector(7 downto 0);
    signal call40_318 : std_logic_vector(7 downto 0);
    signal call42_337 : std_logic_vector(7 downto 0);
    signal call44_356 : std_logic_vector(7 downto 0);
    signal call69_582 : std_logic_vector(7 downto 0);
    signal call72_595 : std_logic_vector(7 downto 0);
    signal call77_613 : std_logic_vector(7 downto 0);
    signal call83_631 : std_logic_vector(7 downto 0);
    signal call89_649 : std_logic_vector(7 downto 0);
    signal call95_667 : std_logic_vector(7 downto 0);
    signal call_37 : std_logic_vector(7 downto 0);
    signal cmp12223_174 : std_logic_vector(0 downto 0);
    signal cmp124208_522 : std_logic_vector(0 downto 0);
    signal cmp12_240 : std_logic_vector(0 downto 0);
    signal cmp191204_998 : std_logic_vector(0 downto 0);
    signal cmp227_58 : std_logic_vector(0 downto 0);
    signal cmp65213_501 : std_logic_vector(0 downto 0);
    signal cmp_130 : std_logic_vector(0 downto 0);
    signal conv103_689 : std_logic_vector(63 downto 0);
    signal conv109_707 : std_logic_vector(63 downto 0);
    signal conv130_796 : std_logic_vector(63 downto 0);
    signal conv135_809 : std_logic_vector(63 downto 0);
    signal conv141_827 : std_logic_vector(63 downto 0);
    signal conv147_845 : std_logic_vector(63 downto 0);
    signal conv153_863 : std_logic_vector(63 downto 0);
    signal conv159_881 : std_logic_vector(63 downto 0);
    signal conv165_899 : std_logic_vector(63 downto 0);
    signal conv16_215 : std_logic_vector(31 downto 0);
    signal conv171_917 : std_logic_vector(63 downto 0);
    signal conv30218_256 : std_logic_vector(15 downto 0);
    signal conv30220_266 : std_logic_vector(15 downto 0);
    signal conv30_288 : std_logic_vector(15 downto 0);
    signal conv30x_xlcssa_308 : std_logic_vector(15 downto 0);
    signal conv41_322 : std_logic_vector(31 downto 0);
    signal conv4229_65 : std_logic_vector(31 downto 0);
    signal conv4231_82 : std_logic_vector(31 downto 0);
    signal conv43_341 : std_logic_vector(31 downto 0);
    signal conv45_360 : std_logic_vector(31 downto 0);
    signal conv4_137 : std_logic_vector(31 downto 0);
    signal conv4x_xlcssa1_145 : std_logic_vector(31 downto 0);
    signal conv4x_xlcssa_152 : std_logic_vector(31 downto 0);
    signal conv51_422 : std_logic_vector(63 downto 0);
    signal conv60_489 : std_logic_vector(63 downto 0);
    signal conv70_586 : std_logic_vector(63 downto 0);
    signal conv74_599 : std_logic_vector(63 downto 0);
    signal conv79_617 : std_logic_vector(63 downto 0);
    signal conv85_635 : std_logic_vector(63 downto 0);
    signal conv91_653 : std_logic_vector(63 downto 0);
    signal conv97_671 : std_logic_vector(63 downto 0);
    signal conv_41 : std_logic_vector(31 downto 0);
    signal exitcond10_727 : std_logic_vector(0 downto 0);
    signal exitcond19_937 : std_logic_vector(0 downto 0);
    signal exitcond20_1073 : std_logic_vector(0 downto 0);
    signal exitcond_300 : std_logic_vector(0 downto 0);
    signal iNsTr_13_121 : std_logic_vector(31 downto 0);
    signal iNsTr_1_47 : std_logic_vector(31 downto 0);
    signal iNsTr_21_231 : std_logic_vector(31 downto 0);
    signal iNsTr_26_330 : std_logic_vector(31 downto 0);
    signal iNsTr_29_349 : std_logic_vector(31 downto 0);
    signal iNsTr_32_368 : std_logic_vector(31 downto 0);
    signal iNsTr_34_380 : std_logic_vector(31 downto 0);
    signal iNsTr_35_392 : std_logic_vector(31 downto 0);
    signal iNsTr_36_404 : std_logic_vector(31 downto 0);
    signal iNsTr_37_430 : std_logic_vector(31 downto 0);
    signal iNsTr_38_442 : std_logic_vector(31 downto 0);
    signal iNsTr_39_454 : std_logic_vector(31 downto 0);
    signal iNsTr_40_466 : std_logic_vector(31 downto 0);
    signal iNsTr_45_954 : std_logic_vector(31 downto 0);
    signal iNsTr_46_966 : std_logic_vector(31 downto 0);
    signal iNsTr_47_978 : std_logic_vector(31 downto 0);
    signal iNsTr_5_164 : std_logic_vector(31 downto 0);
    signal iNsTr_60_1027 : std_logic_vector(63 downto 0);
    signal inc22_201 : std_logic_vector(31 downto 0);
    signal inc_98 : std_logic_vector(31 downto 0);
    signal indvar240_775 : std_logic_vector(63 downto 0);
    signal indvar250_565 : std_logic_vector(63 downto 0);
    signal indvar260_259 : std_logic_vector(63 downto 0);
    signal indvar263_184 : std_logic_vector(63 downto 0);
    signal indvar268_75 : std_logic_vector(63 downto 0);
    signal indvar_1043 : std_logic_vector(63 downto 0);
    signal indvarx_xnext241_932 : std_logic_vector(63 downto 0);
    signal indvarx_xnext251_722 : std_logic_vector(63 downto 0);
    signal indvarx_xnext261_294 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1068 : std_logic_vector(63 downto 0);
    signal mul184_987 : std_logic_vector(31 downto 0);
    signal mul186_992 : std_logic_vector(31 downto 0);
    signal mul50_418 : std_logic_vector(31 downto 0);
    signal mul55_475 : std_logic_vector(31 downto 0);
    signal mul57_480 : std_logic_vector(31 downto 0);
    signal mul59_485 : std_logic_vector(31 downto 0);
    signal mul_413 : std_logic_vector(31 downto 0);
    signal ptr_deref_1059_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1059_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1059_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1059_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1059_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1059_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_107_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_107_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_107_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_107_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_107_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_107_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_124_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_124_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_124_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_124_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_124_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_166_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_166_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_166_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_166_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_166_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_166_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_217_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_217_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_217_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_217_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_217_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_217_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_234_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_234_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_234_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_234_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_234_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_279_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_279_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_279_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_279_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_279_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_279_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_332_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_332_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_332_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_332_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_332_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_332_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_351_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_351_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_351_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_351_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_351_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_351_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_370_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_370_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_370_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_370_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_370_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_370_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_383_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_383_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_383_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_383_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_383_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_395_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_395_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_395_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_395_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_395_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_407_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_407_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_407_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_407_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_407_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_433_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_433_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_433_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_433_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_433_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_445_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_445_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_445_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_445_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_445_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_457_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_457_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_457_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_457_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_457_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_469_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_469_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_469_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_469_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_469_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_49_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_49_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_49_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_49_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_49_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_49_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_714_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_714_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_714_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_714_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_714_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_714_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_924_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_924_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_924_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_924_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_924_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_924_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_957_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_957_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_957_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_957_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_957_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_969_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_969_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_969_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_969_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_969_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_981_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_981_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_981_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_981_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_981_word_offset_0 : std_logic_vector(6 downto 0);
    signal shl100_682 : std_logic_vector(63 downto 0);
    signal shl106_700 : std_logic_vector(63 downto 0);
    signal shl132_802 : std_logic_vector(63 downto 0);
    signal shl138_820 : std_logic_vector(63 downto 0);
    signal shl144_838 : std_logic_vector(63 downto 0);
    signal shl150_856 : std_logic_vector(63 downto 0);
    signal shl156_874 : std_logic_vector(63 downto 0);
    signal shl162_892 : std_logic_vector(63 downto 0);
    signal shl168_910 : std_logic_vector(63 downto 0);
    signal shl76_610 : std_logic_vector(63 downto 0);
    signal shl82_628 : std_logic_vector(63 downto 0);
    signal shl88_646 : std_logic_vector(63 downto 0);
    signal shl94_664 : std_logic_vector(63 downto 0);
    signal shl_592 : std_logic_vector(63 downto 0);
    signal shr123207x_xmask_516 : std_logic_vector(63 downto 0);
    signal shr212x_xmask_495 : std_logic_vector(63 downto 0);
    signal tmp11_235 : std_logic_vector(31 downto 0);
    signal tmp12_739 : std_logic_vector(31 downto 0);
    signal tmp13_744 : std_logic_vector(31 downto 0);
    signal tmp14_749 : std_logic_vector(31 downto 0);
    signal tmp15_753 : std_logic_vector(63 downto 0);
    signal tmp16_759 : std_logic_vector(63 downto 0);
    signal tmp17_765 : std_logic_vector(0 downto 0);
    signal tmp182_958 : std_logic_vector(31 downto 0);
    signal tmp183_970 : std_logic_vector(31 downto 0);
    signal tmp185_982 : std_logic_vector(31 downto 0);
    signal tmp1_125 : std_logic_vector(31 downto 0);
    signal tmp235_1011 : std_logic_vector(31 downto 0);
    signal tmp235x_xop_1023 : std_logic_vector(31 downto 0);
    signal tmp236_1017 : std_logic_vector(0 downto 0);
    signal tmp239_1040 : std_logic_vector(63 downto 0);
    signal tmp265_225 : std_logic_vector(63 downto 0);
    signal tmp270_115 : std_logic_vector(63 downto 0);
    signal tmp3_197 : std_logic_vector(63 downto 0);
    signal tmp47_384 : std_logic_vector(31 downto 0);
    signal tmp48_396 : std_logic_vector(31 downto 0);
    signal tmp49_408 : std_logic_vector(31 downto 0);
    signal tmp53_434 : std_logic_vector(31 downto 0);
    signal tmp54_446 : std_logic_vector(31 downto 0);
    signal tmp56_458 : std_logic_vector(31 downto 0);
    signal tmp58_470 : std_logic_vector(31 downto 0);
    signal tmp5_534 : std_logic_vector(31 downto 0);
    signal tmp6_539 : std_logic_vector(31 downto 0);
    signal tmp7_543 : std_logic_vector(63 downto 0);
    signal tmp8_549 : std_logic_vector(63 downto 0);
    signal tmp9_555 : std_logic_vector(0 downto 0);
    signal tmp_94 : std_logic_vector(63 downto 0);
    signal type_cast_1009_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1015_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1021_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1031_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1038_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1047_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1049_wire : std_logic_vector(63 downto 0);
    signal type_cast_1061_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1066_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_113_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_148_wire : std_logic_vector(31 downto 0);
    signal type_cast_155_wire : std_logic_vector(31 downto 0);
    signal type_cast_157_wire : std_logic_vector(31 downto 0);
    signal type_cast_172_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_187_wire : std_logic_vector(63 downto 0);
    signal type_cast_190_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_195_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_223_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_263_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_265_wire : std_logic_vector(63 downto 0);
    signal type_cast_269_wire : std_logic_vector(15 downto 0);
    signal type_cast_271_wire : std_logic_vector(15 downto 0);
    signal type_cast_292_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_298_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_311_wire : std_logic_vector(15 downto 0);
    signal type_cast_493_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_514_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_547_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_55_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_560_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_569_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_571_wire : std_logic_vector(63 downto 0);
    signal type_cast_590_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_608_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_644_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_662_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_680_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_698_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_720_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_757_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_763_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_770_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_779_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_781_wire : std_logic_vector(63 downto 0);
    signal type_cast_78_wire : std_logic_vector(63 downto 0);
    signal type_cast_800_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_818_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_81_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_836_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_854_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_85_wire : std_logic_vector(31 downto 0);
    signal type_cast_872_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_87_wire : std_logic_vector(31 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_92_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_930_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_996_wire_constant : std_logic_vector(31 downto 0);
    signal umax18_772 : std_logic_vector(63 downto 0);
    signal umax_562 : std_logic_vector(63 downto 0);
    signal xx_xop_1033 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_padding_313_word_address_0 <= "0";
    array_obj_ref_103_constant_part_of_offset <= "0000010";
    array_obj_ref_103_offset_scale_factor_0 <= "1000000";
    array_obj_ref_103_offset_scale_factor_1 <= "0000001";
    array_obj_ref_103_resized_base_address <= "0000000";
    array_obj_ref_1055_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1055_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1055_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1055_resized_base_address <= "00000000000000";
    array_obj_ref_206_constant_part_of_offset <= "0000010";
    array_obj_ref_206_offset_scale_factor_0 <= "1000000";
    array_obj_ref_206_offset_scale_factor_1 <= "0000001";
    array_obj_ref_206_resized_base_address <= "0000000";
    array_obj_ref_275_offset_scale_factor_0 <= "1";
    array_obj_ref_275_resized_base_address <= "0";
    array_obj_ref_577_constant_part_of_offset <= "00000000000000";
    array_obj_ref_577_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_577_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_577_resized_base_address <= "00000000000000";
    array_obj_ref_787_constant_part_of_offset <= "00000100001";
    array_obj_ref_787_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_787_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_787_resized_base_address <= "00000000000";
    iNsTr_13_121 <= "00000000000000000000000000000001";
    iNsTr_1_47 <= "00000000000000000000000000000001";
    iNsTr_21_231 <= "00000000000000000000000000000001";
    iNsTr_26_330 <= "00000000000000000000000000000010";
    iNsTr_29_349 <= "00000000000000000000000000000011";
    iNsTr_32_368 <= "00000000000000000000000000000100";
    iNsTr_34_380 <= "00000000000000000000000000000010";
    iNsTr_35_392 <= "00000000000000000000000000000011";
    iNsTr_36_404 <= "00000000000000000000000000000100";
    iNsTr_37_430 <= "00000000000000000000000000000010";
    iNsTr_38_442 <= "00000000000000000000000000000011";
    iNsTr_39_454 <= "00000000000000000000000000000100";
    iNsTr_40_466 <= "00000000000000000000000000000101";
    iNsTr_45_954 <= "00000000000000000000000000000010";
    iNsTr_46_966 <= "00000000000000000000000000000011";
    iNsTr_47_978 <= "00000000000000000000000000000100";
    iNsTr_5_164 <= "00000000000000000000000000000001";
    ptr_deref_1059_word_offset_0 <= "00000000000000";
    ptr_deref_107_word_offset_0 <= "0000000";
    ptr_deref_124_word_offset_0 <= "0000000";
    ptr_deref_166_word_offset_0 <= "0000000";
    ptr_deref_217_word_offset_0 <= "0000000";
    ptr_deref_234_word_offset_0 <= "0000000";
    ptr_deref_279_word_offset_0 <= "0";
    ptr_deref_332_word_offset_0 <= "0000000";
    ptr_deref_351_word_offset_0 <= "0000000";
    ptr_deref_370_word_offset_0 <= "0000000";
    ptr_deref_383_word_offset_0 <= "0000000";
    ptr_deref_395_word_offset_0 <= "0000000";
    ptr_deref_407_word_offset_0 <= "0000000";
    ptr_deref_433_word_offset_0 <= "0000000";
    ptr_deref_445_word_offset_0 <= "0000000";
    ptr_deref_457_word_offset_0 <= "0000000";
    ptr_deref_469_word_offset_0 <= "0000000";
    ptr_deref_49_word_offset_0 <= "0000000";
    ptr_deref_714_word_offset_0 <= "00000000000000";
    ptr_deref_924_word_offset_0 <= "00000000000";
    ptr_deref_957_word_offset_0 <= "0000000";
    ptr_deref_969_word_offset_0 <= "0000000";
    ptr_deref_981_word_offset_0 <= "0000000";
    type_cast_1009_wire_constant <= "00000000000000000000000000000010";
    type_cast_1015_wire_constant <= "00000000000000000000000000000001";
    type_cast_1021_wire_constant <= "11111111111111111111111111111111";
    type_cast_1031_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1038_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1047_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1061_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1066_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_113_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_172_wire_constant <= "00000000000000000000000000000000";
    type_cast_190_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_195_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_223_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_263_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_292_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_298_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_493_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_499_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_514_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_520_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_547_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_553_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_55_wire_constant <= "00000000";
    type_cast_560_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_569_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_590_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_608_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_626_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_644_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_662_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_680_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_698_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_720_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_757_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_763_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_770_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_779_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_800_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_818_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_81_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_836_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_854_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_872_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_890_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_92_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_930_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_996_wire_constant <= "00000000000000000000000000000011";
    phi_stmt_1043: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1047_wire_constant & type_cast_1049_wire;
      req <= phi_stmt_1043_req_0 & phi_stmt_1043_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1043",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1043_ack_0,
          idata => idata,
          odata => indvar_1043,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1043
    phi_stmt_145: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_148_wire;
      req(0) <= phi_stmt_145_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_145",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_145_ack_0,
          idata => idata,
          odata => conv4x_xlcssa1_145,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_145
    phi_stmt_152: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_155_wire & type_cast_157_wire;
      req <= phi_stmt_152_req_0 & phi_stmt_152_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_152",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_152_ack_0,
          idata => idata,
          odata => conv4x_xlcssa_152,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_152
    phi_stmt_184: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_187_wire & type_cast_190_wire_constant;
      req <= phi_stmt_184_req_0 & phi_stmt_184_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_184",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_184_ack_0,
          idata => idata,
          odata => indvar263_184,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_184
    phi_stmt_259: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_263_wire_constant & type_cast_265_wire;
      req <= phi_stmt_259_req_0 & phi_stmt_259_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_259",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_259_ack_0,
          idata => idata,
          odata => indvar260_259,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_259
    phi_stmt_266: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_269_wire & type_cast_271_wire;
      req <= phi_stmt_266_req_0 & phi_stmt_266_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_266",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_266_ack_0,
          idata => idata,
          odata => conv30220_266,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_266
    phi_stmt_308: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_311_wire;
      req(0) <= phi_stmt_308_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_308",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_308_ack_0,
          idata => idata,
          odata => conv30x_xlcssa_308,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_308
    phi_stmt_565: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_569_wire_constant & type_cast_571_wire;
      req <= phi_stmt_565_req_0 & phi_stmt_565_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_565",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_565_ack_0,
          idata => idata,
          odata => indvar250_565,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_565
    phi_stmt_75: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_78_wire & type_cast_81_wire_constant;
      req <= phi_stmt_75_req_0 & phi_stmt_75_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_75",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_75_ack_0,
          idata => idata,
          odata => indvar268_75,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_75
    phi_stmt_775: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_779_wire_constant & type_cast_781_wire;
      req <= phi_stmt_775_req_0 & phi_stmt_775_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_775",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_775_ack_0,
          idata => idata,
          odata => indvar240_775,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_775
    phi_stmt_82: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_85_wire & type_cast_87_wire;
      req <= phi_stmt_82_req_0 & phi_stmt_82_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_82",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_82_ack_0,
          idata => idata,
          odata => conv4231_82,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_82
    -- flow-through select operator MUX_1039_inst
    tmp239_1040 <= xx_xop_1033 when (tmp236_1017(0) /=  '0') else type_cast_1038_wire_constant;
    -- flow-through select operator MUX_561_inst
    umax_562 <= tmp8_549 when (tmp9_555(0) /=  '0') else type_cast_560_wire_constant;
    -- flow-through select operator MUX_771_inst
    umax18_772 <= tmp16_759 when (tmp17_765(0) /=  '0') else type_cast_770_wire_constant;
    addr_of_104_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_104_final_reg_req_0;
      addr_of_104_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_104_final_reg_req_1;
      addr_of_104_final_reg_ack_1<= rack(0);
      addr_of_104_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_104_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_103_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1056_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1056_final_reg_req_0;
      addr_of_1056_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1056_final_reg_req_1;
      addr_of_1056_final_reg_ack_1<= rack(0);
      addr_of_1056_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1056_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1055_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx196_1057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_207_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_207_final_reg_req_0;
      addr_of_207_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_207_final_reg_req_1;
      addr_of_207_final_reg_ack_1<= rack(0);
      addr_of_207_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_207_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_206_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx19_208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_276_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_276_final_reg_req_0;
      addr_of_276_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_276_final_reg_req_1;
      addr_of_276_final_reg_ack_1<= rack(0);
      addr_of_276_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_276_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_275_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx33_277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_578_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_578_final_reg_req_0;
      addr_of_578_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_578_final_reg_req_1;
      addr_of_578_final_reg_ack_1<= rack(0);
      addr_of_578_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_578_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_577_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx114_579,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_788_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_788_final_reg_req_0;
      addr_of_788_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_788_final_reg_req_1;
      addr_of_788_final_reg_ack_1<= rack(0);
      addr_of_788_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_788_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_787_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx176_789,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1026_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1026_inst_req_0;
      type_cast_1026_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1026_inst_req_1;
      type_cast_1026_inst_ack_1<= rack(0);
      type_cast_1026_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1026_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp235x_xop_1023,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_60_1027,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1049_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1049_inst_req_0;
      type_cast_1049_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1049_inst_req_1;
      type_cast_1049_inst_ack_1<= rack(0);
      type_cast_1049_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1049_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1068,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1049_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1085_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1085_inst_req_0;
      type_cast_1085_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1085_inst_req_1;
      type_cast_1085_inst_ack_1<= rack(0);
      type_cast_1085_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1085_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul50_418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_136_inst_req_0;
      type_cast_136_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_136_inst_req_1;
      type_cast_136_inst_ack_1<= rack(0);
      type_cast_136_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_136_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_137,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_148_inst_req_0;
      type_cast_148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_148_inst_req_1;
      type_cast_148_inst_ack_1<= rack(0);
      type_cast_148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_148_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_155_inst_req_0;
      type_cast_155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_155_inst_req_1;
      type_cast_155_inst_ack_1<= rack(0);
      type_cast_155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4229_65,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_155_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_157_inst_req_0;
      type_cast_157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_157_inst_req_1;
      type_cast_157_inst_ack_1<= rack(0);
      type_cast_157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4x_xlcssa1_145,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_157_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_187_inst_req_0;
      type_cast_187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_187_inst_req_1;
      type_cast_187_inst_ack_1<= rack(0);
      type_cast_187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp265_225,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_187_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_200_inst_req_0;
      type_cast_200_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_200_inst_req_1;
      type_cast_200_inst_ack_1<= rack(0);
      type_cast_200_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_200_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_197,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc22_201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_214_inst_req_0;
      type_cast_214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_214_inst_req_1;
      type_cast_214_inst_ack_1<= rack(0);
      type_cast_214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_255_inst_req_0;
      type_cast_255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_255_inst_req_1;
      type_cast_255_inst_ack_1<= rack(0);
      type_cast_255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29217_252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30218_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_265_inst_req_0;
      type_cast_265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_265_inst_req_1;
      type_cast_265_inst_ack_1<= rack(0);
      type_cast_265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext261_294,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_265_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_269_inst_req_0;
      type_cast_269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_269_inst_req_1;
      type_cast_269_inst_ack_1<= rack(0);
      type_cast_269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30218_256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_269_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_271_inst_req_0;
      type_cast_271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_271_inst_req_1;
      type_cast_271_inst_ack_1<= rack(0);
      type_cast_271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_271_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_271_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_287_inst_req_0;
      type_cast_287_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_287_inst_req_1;
      type_cast_287_inst_ack_1<= rack(0);
      type_cast_287_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_287_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29_284,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_311_inst_req_0;
      type_cast_311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_311_inst_req_1;
      type_cast_311_inst_ack_1<= rack(0);
      type_cast_311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_311_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_321_inst_req_0;
      type_cast_321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_321_inst_req_1;
      type_cast_321_inst_ack_1<= rack(0);
      type_cast_321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call40_318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_340_inst_req_0;
      type_cast_340_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_340_inst_req_1;
      type_cast_340_inst_ack_1<= rack(0);
      type_cast_340_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_340_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_341,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_359_inst_req_0;
      type_cast_359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_359_inst_req_1;
      type_cast_359_inst_ack_1<= rack(0);
      type_cast_359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_360,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_40_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_40_inst_req_0;
      type_cast_40_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_40_inst_req_1;
      type_cast_40_inst_ack_1<= rack(0);
      type_cast_40_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_40_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_37,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_41,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_421_inst_req_0;
      type_cast_421_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_421_inst_req_1;
      type_cast_421_inst_ack_1<= rack(0);
      type_cast_421_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_421_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul50_418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_488_inst_req_0;
      type_cast_488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_488_inst_req_1;
      type_cast_488_inst_ack_1<= rack(0);
      type_cast_488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul59_485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_542_inst_req_0;
      type_cast_542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_542_inst_req_1;
      type_cast_542_inst_ack_1<= rack(0);
      type_cast_542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_542_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp6_539,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp7_543,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_571_inst_req_0;
      type_cast_571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_571_inst_req_1;
      type_cast_571_inst_ack_1<= rack(0);
      type_cast_571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_571_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext251_722,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_571_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_585_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_585_inst_req_0;
      type_cast_585_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_585_inst_req_1;
      type_cast_585_inst_ack_1<= rack(0);
      type_cast_585_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_585_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call69_582,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_586,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_598_inst_req_0;
      type_cast_598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_598_inst_req_1;
      type_cast_598_inst_ack_1<= rack(0);
      type_cast_598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call72_595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_616_inst_req_0;
      type_cast_616_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_616_inst_req_1;
      type_cast_616_inst_ack_1<= rack(0);
      type_cast_616_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_616_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call77_613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_617,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_634_inst_req_0;
      type_cast_634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_634_inst_req_1;
      type_cast_634_inst_ack_1<= rack(0);
      type_cast_634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call83_631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3228_61,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4229_65,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_652_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_652_inst_req_0;
      type_cast_652_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_652_inst_req_1;
      type_cast_652_inst_ack_1<= rack(0);
      type_cast_652_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_652_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_653,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_670_inst_req_0;
      type_cast_670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_670_inst_req_1;
      type_cast_670_inst_ack_1<= rack(0);
      type_cast_670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_667,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_688_inst_req_0;
      type_cast_688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_688_inst_req_1;
      type_cast_688_inst_ack_1<= rack(0);
      type_cast_688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_685,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_706_inst_req_0;
      type_cast_706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_706_inst_req_1;
      type_cast_706_inst_ack_1<= rack(0);
      type_cast_706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_707,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_752_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_752_inst_req_0;
      type_cast_752_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_752_inst_req_1;
      type_cast_752_inst_ack_1<= rack(0);
      type_cast_752_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_752_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_749,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_753,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_781_inst_req_0;
      type_cast_781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_781_inst_req_1;
      type_cast_781_inst_ack_1<= rack(0);
      type_cast_781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext241_932,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_781_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_78_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_78_inst_req_0;
      type_cast_78_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_78_inst_req_1;
      type_cast_78_inst_ack_1<= rack(0);
      type_cast_78_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_78_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp270_115,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_78_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_795_inst_req_0;
      type_cast_795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_795_inst_req_1;
      type_cast_795_inst_ack_1<= rack(0);
      type_cast_795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_808_inst_req_0;
      type_cast_808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_808_inst_req_1;
      type_cast_808_inst_ack_1<= rack(0);
      type_cast_808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_805,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_809,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_826_inst_req_0;
      type_cast_826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_826_inst_req_1;
      type_cast_826_inst_ack_1<= rack(0);
      type_cast_826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call139_823,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_827,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_844_inst_req_0;
      type_cast_844_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_844_inst_req_1;
      type_cast_844_inst_ack_1<= rack(0);
      type_cast_844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_841,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_845,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_85_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_85_inst_req_0;
      type_cast_85_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_85_inst_req_1;
      type_cast_85_inst_ack_1<= rack(0);
      type_cast_85_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_85_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_85_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_862_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_862_inst_req_0;
      type_cast_862_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_862_inst_req_1;
      type_cast_862_inst_ack_1<= rack(0);
      type_cast_862_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_862_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call151_859,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_863,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_87_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_87_inst_req_0;
      type_cast_87_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_87_inst_req_1;
      type_cast_87_inst_ack_1<= rack(0);
      type_cast_87_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_87_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4229_65,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_87_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_880_inst_req_0;
      type_cast_880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_880_inst_req_1;
      type_cast_880_inst_ack_1<= rack(0);
      type_cast_880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call157_877,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_898_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_898_inst_req_0;
      type_cast_898_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_898_inst_req_1;
      type_cast_898_inst_ack_1<= rack(0);
      type_cast_898_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_898_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call163_895,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_899,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_916_inst_req_0;
      type_cast_916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_916_inst_req_1;
      type_cast_916_inst_ack_1<= rack(0);
      type_cast_916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_917,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_97_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_97_inst_req_0;
      type_cast_97_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_97_inst_req_1;
      type_cast_97_inst_ack_1<= rack(0);
      type_cast_97_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_97_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_94,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_98,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_padding_313_gather_scatter
    process(conv30x_xlcssa_308) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv30x_xlcssa_308;
      ov(15 downto 0) := iv;
      STORE_padding_313_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_103_index_1_rename
    process(R_indvar268_102_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar268_102_resized;
      ov(6 downto 0) := iv;
      R_indvar268_102_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_103_index_1_resize
    process(indvar268_75) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar268_75;
      ov := iv(6 downto 0);
      R_indvar268_102_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_103_root_address_inst
    process(array_obj_ref_103_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_103_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_103_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1055_index_1_rename
    process(R_indvar_1054_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1054_resized;
      ov(13 downto 0) := iv;
      R_indvar_1054_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1055_index_1_resize
    process(indvar_1043) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1043;
      ov := iv(13 downto 0);
      R_indvar_1054_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1055_root_address_inst
    process(array_obj_ref_1055_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1055_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1055_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_206_index_1_rename
    process(R_indvar263_205_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar263_205_resized;
      ov(6 downto 0) := iv;
      R_indvar263_205_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_206_index_1_resize
    process(indvar263_184) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar263_184;
      ov := iv(6 downto 0);
      R_indvar263_205_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_206_root_address_inst
    process(array_obj_ref_206_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_206_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_206_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_275_index_0_rename
    process(R_indvar260_274_resized) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar260_274_resized;
      ov(0 downto 0) := iv;
      R_indvar260_274_scaled <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_275_index_0_resize
    process(indvar260_259) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar260_259;
      ov := iv(0 downto 0);
      R_indvar260_274_resized <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_275_index_offset
    process(R_indvar260_274_scaled) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar260_274_scaled;
      ov(0 downto 0) := iv;
      array_obj_ref_275_final_offset <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_275_root_address_inst
    process(array_obj_ref_275_final_offset) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_275_final_offset;
      ov(0 downto 0) := iv;
      array_obj_ref_275_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_577_index_1_rename
    process(R_indvar250_576_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar250_576_resized;
      ov(13 downto 0) := iv;
      R_indvar250_576_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_577_index_1_resize
    process(indvar250_565) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar250_565;
      ov := iv(13 downto 0);
      R_indvar250_576_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_577_root_address_inst
    process(array_obj_ref_577_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_577_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_577_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_787_index_1_rename
    process(R_indvar240_786_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar240_786_resized;
      ov(10 downto 0) := iv;
      R_indvar240_786_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_787_index_1_resize
    process(indvar240_775) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar240_775;
      ov := iv(10 downto 0);
      R_indvar240_786_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_787_root_address_inst
    process(array_obj_ref_787_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_787_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_787_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1059_addr_0
    process(ptr_deref_1059_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1059_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1059_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1059_base_resize
    process(arrayidx196_1057) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx196_1057;
      ov := iv(13 downto 0);
      ptr_deref_1059_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1059_gather_scatter
    process(type_cast_1061_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1061_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1059_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1059_root_address_inst
    process(ptr_deref_1059_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1059_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1059_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_107_addr_0
    process(ptr_deref_107_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_107_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_107_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_107_base_resize
    process(arrayidx_105) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_105;
      ov := iv(6 downto 0);
      ptr_deref_107_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_107_gather_scatter
    process(conv4231_82) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4231_82;
      ov(31 downto 0) := iv;
      ptr_deref_107_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_107_root_address_inst
    process(ptr_deref_107_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_107_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_107_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_124_addr_0
    process(ptr_deref_124_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_124_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_124_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_124_base_resize
    process(iNsTr_13_121) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_13_121;
      ov := iv(6 downto 0);
      ptr_deref_124_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_124_gather_scatter
    process(ptr_deref_124_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_124_data_0;
      ov(31 downto 0) := iv;
      tmp1_125 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_124_root_address_inst
    process(ptr_deref_124_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_124_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_124_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_166_addr_0
    process(ptr_deref_166_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_166_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_166_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_166_base_resize
    process(iNsTr_5_164) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_164;
      ov := iv(6 downto 0);
      ptr_deref_166_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_166_gather_scatter
    process(conv4x_xlcssa_152) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4x_xlcssa_152;
      ov(31 downto 0) := iv;
      ptr_deref_166_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_166_root_address_inst
    process(ptr_deref_166_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_166_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_166_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_217_addr_0
    process(ptr_deref_217_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_217_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_217_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_217_base_resize
    process(arrayidx19_208) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx19_208;
      ov := iv(6 downto 0);
      ptr_deref_217_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_217_gather_scatter
    process(conv16_215) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv16_215;
      ov(31 downto 0) := iv;
      ptr_deref_217_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_217_root_address_inst
    process(ptr_deref_217_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_217_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_217_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_234_addr_0
    process(ptr_deref_234_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_234_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_234_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_234_base_resize
    process(iNsTr_21_231) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_231;
      ov := iv(6 downto 0);
      ptr_deref_234_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_234_gather_scatter
    process(ptr_deref_234_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_234_data_0;
      ov(31 downto 0) := iv;
      tmp11_235 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_234_root_address_inst
    process(ptr_deref_234_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_234_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_234_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_279_addr_0
    process(ptr_deref_279_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_279_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_279_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_279_base_resize
    process(arrayidx33_277) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx33_277;
      ov := iv(0 downto 0);
      ptr_deref_279_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_279_gather_scatter
    process(conv30220_266) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv30220_266;
      ov(15 downto 0) := iv;
      ptr_deref_279_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_279_root_address_inst
    process(ptr_deref_279_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_279_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_279_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_332_addr_0
    process(ptr_deref_332_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_332_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_332_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_332_base_resize
    process(iNsTr_26_330) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_330;
      ov := iv(6 downto 0);
      ptr_deref_332_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_332_gather_scatter
    process(conv41_322) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv41_322;
      ov(31 downto 0) := iv;
      ptr_deref_332_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_332_root_address_inst
    process(ptr_deref_332_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_332_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_332_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_351_addr_0
    process(ptr_deref_351_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_351_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_351_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_351_base_resize
    process(iNsTr_29_349) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_29_349;
      ov := iv(6 downto 0);
      ptr_deref_351_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_351_gather_scatter
    process(conv43_341) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv43_341;
      ov(31 downto 0) := iv;
      ptr_deref_351_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_351_root_address_inst
    process(ptr_deref_351_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_351_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_351_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_370_addr_0
    process(ptr_deref_370_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_370_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_370_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_370_base_resize
    process(iNsTr_32_368) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_32_368;
      ov := iv(6 downto 0);
      ptr_deref_370_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_370_gather_scatter
    process(conv45_360) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv45_360;
      ov(31 downto 0) := iv;
      ptr_deref_370_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_370_root_address_inst
    process(ptr_deref_370_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_370_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_370_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_addr_0
    process(ptr_deref_383_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_383_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_383_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_base_resize
    process(iNsTr_34_380) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_380;
      ov := iv(6 downto 0);
      ptr_deref_383_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_gather_scatter
    process(ptr_deref_383_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_383_data_0;
      ov(31 downto 0) := iv;
      tmp47_384 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_root_address_inst
    process(ptr_deref_383_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_383_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_383_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_395_addr_0
    process(ptr_deref_395_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_395_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_395_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_395_base_resize
    process(iNsTr_35_392) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_35_392;
      ov := iv(6 downto 0);
      ptr_deref_395_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_395_gather_scatter
    process(ptr_deref_395_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_395_data_0;
      ov(31 downto 0) := iv;
      tmp48_396 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_395_root_address_inst
    process(ptr_deref_395_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_395_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_395_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_addr_0
    process(ptr_deref_407_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_407_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_base_resize
    process(iNsTr_36_404) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_36_404;
      ov := iv(6 downto 0);
      ptr_deref_407_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_gather_scatter
    process(ptr_deref_407_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_data_0;
      ov(31 downto 0) := iv;
      tmp49_408 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_root_address_inst
    process(ptr_deref_407_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_407_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_433_addr_0
    process(ptr_deref_433_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_433_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_433_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_433_base_resize
    process(iNsTr_37_430) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_430;
      ov := iv(6 downto 0);
      ptr_deref_433_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_433_gather_scatter
    process(ptr_deref_433_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_433_data_0;
      ov(31 downto 0) := iv;
      tmp53_434 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_433_root_address_inst
    process(ptr_deref_433_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_433_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_433_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_445_addr_0
    process(ptr_deref_445_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_445_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_445_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_445_base_resize
    process(iNsTr_38_442) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_442;
      ov := iv(6 downto 0);
      ptr_deref_445_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_445_gather_scatter
    process(ptr_deref_445_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_445_data_0;
      ov(31 downto 0) := iv;
      tmp54_446 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_445_root_address_inst
    process(ptr_deref_445_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_445_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_445_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_457_addr_0
    process(ptr_deref_457_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_457_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_457_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_457_base_resize
    process(iNsTr_39_454) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_39_454;
      ov := iv(6 downto 0);
      ptr_deref_457_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_457_gather_scatter
    process(ptr_deref_457_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_457_data_0;
      ov(31 downto 0) := iv;
      tmp56_458 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_457_root_address_inst
    process(ptr_deref_457_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_457_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_457_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_469_addr_0
    process(ptr_deref_469_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_469_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_469_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_469_base_resize
    process(iNsTr_40_466) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_466;
      ov := iv(6 downto 0);
      ptr_deref_469_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_469_gather_scatter
    process(ptr_deref_469_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_469_data_0;
      ov(31 downto 0) := iv;
      tmp58_470 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_469_root_address_inst
    process(ptr_deref_469_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_469_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_469_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_addr_0
    process(ptr_deref_49_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_49_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_49_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_base_resize
    process(iNsTr_1_47) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_47;
      ov := iv(6 downto 0);
      ptr_deref_49_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_gather_scatter
    process(conv_41) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_41;
      ov(31 downto 0) := iv;
      ptr_deref_49_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_root_address_inst
    process(ptr_deref_49_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_49_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_49_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_714_addr_0
    process(ptr_deref_714_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_714_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_714_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_714_base_resize
    process(arrayidx114_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx114_579;
      ov := iv(13 downto 0);
      ptr_deref_714_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_714_gather_scatter
    process(add110_712) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add110_712;
      ov(63 downto 0) := iv;
      ptr_deref_714_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_714_root_address_inst
    process(ptr_deref_714_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_714_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_714_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_924_addr_0
    process(ptr_deref_924_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_924_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_924_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_924_base_resize
    process(arrayidx176_789) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx176_789;
      ov := iv(10 downto 0);
      ptr_deref_924_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_924_gather_scatter
    process(add172_922) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add172_922;
      ov(63 downto 0) := iv;
      ptr_deref_924_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_924_root_address_inst
    process(ptr_deref_924_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_924_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_924_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_957_addr_0
    process(ptr_deref_957_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_957_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_957_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_957_base_resize
    process(iNsTr_45_954) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_45_954;
      ov := iv(6 downto 0);
      ptr_deref_957_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_957_gather_scatter
    process(ptr_deref_957_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_957_data_0;
      ov(31 downto 0) := iv;
      tmp182_958 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_957_root_address_inst
    process(ptr_deref_957_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_957_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_957_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_969_addr_0
    process(ptr_deref_969_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_969_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_969_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_969_base_resize
    process(iNsTr_46_966) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_46_966;
      ov := iv(6 downto 0);
      ptr_deref_969_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_969_gather_scatter
    process(ptr_deref_969_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_969_data_0;
      ov(31 downto 0) := iv;
      tmp183_970 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_969_root_address_inst
    process(ptr_deref_969_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_969_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_969_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_981_addr_0
    process(ptr_deref_981_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_981_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_981_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_981_base_resize
    process(iNsTr_47_978) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_47_978;
      ov := iv(6 downto 0);
      ptr_deref_981_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_981_gather_scatter
    process(ptr_deref_981_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_981_data_0;
      ov(31 downto 0) := iv;
      tmp185_982 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_981_root_address_inst
    process(ptr_deref_981_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_981_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_981_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1074_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond20_1073;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1074_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1074_branch_req_0,
          ack0 => if_stmt_1074_branch_ack_0,
          ack1 => if_stmt_1074_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_138_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_130;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_138_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_138_branch_req_0,
          ack0 => if_stmt_138_branch_ack_0,
          ack1 => if_stmt_138_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_175_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp12223_174;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_175_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_175_branch_req_0,
          ack0 => if_stmt_175_branch_ack_0,
          ack1 => if_stmt_175_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_241_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp12_240;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_241_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_241_branch_req_0,
          ack0 => if_stmt_241_branch_ack_0,
          ack1 => if_stmt_241_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_301_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_300;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_301_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_301_branch_req_0,
          ack0 => if_stmt_301_branch_ack_0,
          ack1 => if_stmt_301_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_502_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp65213_501;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_502_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_502_branch_req_0,
          ack0 => if_stmt_502_branch_ack_0,
          ack1 => if_stmt_502_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_523_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp124208_522;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_523_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_523_branch_req_0,
          ack0 => if_stmt_523_branch_ack_0,
          ack1 => if_stmt_523_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_66_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp227_58;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_66_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_66_branch_req_0,
          ack0 => if_stmt_66_branch_ack_0,
          ack1 => if_stmt_66_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_728_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond10_727;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_728_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_728_branch_req_0,
          ack0 => if_stmt_728_branch_ack_0,
          ack1 => if_stmt_728_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_938_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond19_937;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_938_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_938_branch_req_0,
          ack0 => if_stmt_938_branch_ack_0,
          ack1 => if_stmt_938_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_999_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp191204_998;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_999_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_999_branch_req_0,
          ack0 => if_stmt_999_branch_ack_0,
          ack1 => if_stmt_999_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1022_inst
    process(tmp235_1011) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp235_1011, type_cast_1021_wire_constant, tmp_var);
      tmp235x_xop_1023 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1032_inst
    process(iNsTr_60_1027) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_60_1027, type_cast_1031_wire_constant, tmp_var);
      xx_xop_1033 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1067_inst
    process(indvar_1043) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1043, type_cast_1066_wire_constant, tmp_var);
      indvarx_xnext_1068 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_114_inst
    process(indvar268_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar268_75, type_cast_113_wire_constant, tmp_var);
      tmp270_115 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_196_inst
    process(indvar263_184) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar263_184, type_cast_195_wire_constant, tmp_var);
      tmp3_197 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_224_inst
    process(indvar263_184) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar263_184, type_cast_223_wire_constant, tmp_var);
      tmp265_225 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_293_inst
    process(indvar260_259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar260_259, type_cast_292_wire_constant, tmp_var);
      indvarx_xnext261_294 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_721_inst
    process(indvar250_565) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar250_565, type_cast_720_wire_constant, tmp_var);
      indvarx_xnext251_722 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_931_inst
    process(indvar240_775) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar240_775, type_cast_930_wire_constant, tmp_var);
      indvarx_xnext241_932 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_93_inst
    process(indvar268_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar268_75, type_cast_92_wire_constant, tmp_var);
      tmp_94 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_494_inst
    process(conv51_422) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv51_422, type_cast_493_wire_constant, tmp_var);
      shr212x_xmask_495 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_515_inst
    process(conv60_489) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv60_489, type_cast_514_wire_constant, tmp_var);
      shr123207x_xmask_516 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_173_inst
    process(conv4x_xlcssa_152) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv4x_xlcssa_152, type_cast_172_wire_constant, tmp_var);
      cmp12223_174 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1072_inst
    process(indvarx_xnext_1068, tmp239_1040) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1068, tmp239_1040, tmp_var);
      exitcond20_1073 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_299_inst
    process(indvarx_xnext261_294) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext261_294, type_cast_298_wire_constant, tmp_var);
      exitcond_300 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_500_inst
    process(shr212x_xmask_495) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr212x_xmask_495, type_cast_499_wire_constant, tmp_var);
      cmp65213_501 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_521_inst
    process(shr123207x_xmask_516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr123207x_xmask_516, type_cast_520_wire_constant, tmp_var);
      cmp124208_522 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_726_inst
    process(indvarx_xnext251_722, umax_562) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext251_722, umax_562, tmp_var);
      exitcond10_727 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_936_inst
    process(indvarx_xnext241_932, umax18_772) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext241_932, umax18_772, tmp_var);
      exitcond19_937 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_56_inst
    process(call_37) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(call_37, type_cast_55_wire_constant, tmp_var);
      cmp227_58 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1010_inst
    process(mul186_992) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul186_992, type_cast_1009_wire_constant, tmp_var);
      tmp235_1011 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_548_inst
    process(tmp7_543) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp7_543, type_cast_547_wire_constant, tmp_var);
      tmp8_549 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_758_inst
    process(tmp15_753) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp15_753, type_cast_757_wire_constant, tmp_var);
      tmp16_759 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_412_inst
    process(tmp48_396, tmp47_384) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_396, tmp47_384, tmp_var);
      mul_413 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_417_inst
    process(mul_413, tmp49_408) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_413, tmp49_408, tmp_var);
      mul50_418 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_474_inst
    process(tmp54_446, tmp53_434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_446, tmp53_434, tmp_var);
      mul55_475 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_479_inst
    process(mul55_475, tmp56_458) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul55_475, tmp56_458, tmp_var);
      mul57_480 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_484_inst
    process(mul57_480, tmp58_470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul57_480, tmp58_470, tmp_var);
      mul59_485 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_533_inst
    process(tmp48_396, tmp47_384) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_396, tmp47_384, tmp_var);
      tmp5_534 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_538_inst
    process(tmp5_534, tmp49_408) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp5_534, tmp49_408, tmp_var);
      tmp6_539 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_738_inst
    process(tmp54_446, tmp53_434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_446, tmp53_434, tmp_var);
      tmp12_739 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_743_inst
    process(tmp12_739, tmp56_458) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_739, tmp56_458, tmp_var);
      tmp13_744 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_748_inst
    process(tmp13_744, tmp58_470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_744, tmp58_470, tmp_var);
      tmp14_749 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_986_inst
    process(tmp183_970, tmp182_958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp183_970, tmp182_958, tmp_var);
      mul184_987 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_991_inst
    process(mul184_987, tmp185_982) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul184_987, tmp185_982, tmp_var);
      mul186_992 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_603_inst
    process(shl_592, conv74_599) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_592, conv74_599, tmp_var);
      add_604 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_621_inst
    process(shl76_610, conv79_617) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl76_610, conv79_617, tmp_var);
      add80_622 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_639_inst
    process(shl82_628, conv85_635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl82_628, conv85_635, tmp_var);
      add86_640 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_657_inst
    process(shl88_646, conv91_653) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl88_646, conv91_653, tmp_var);
      add92_658 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_675_inst
    process(shl94_664, conv97_671) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl94_664, conv97_671, tmp_var);
      add98_676 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_693_inst
    process(shl100_682, conv103_689) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_682, conv103_689, tmp_var);
      add104_694 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_711_inst
    process(shl106_700, conv109_707) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl106_700, conv109_707, tmp_var);
      add110_712 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_813_inst
    process(shl132_802, conv135_809) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_802, conv135_809, tmp_var);
      add136_814 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_831_inst
    process(shl138_820, conv141_827) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl138_820, conv141_827, tmp_var);
      add142_832 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_849_inst
    process(shl144_838, conv147_845) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_838, conv147_845, tmp_var);
      add148_850 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_867_inst
    process(shl150_856, conv153_863) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl150_856, conv153_863, tmp_var);
      add154_868 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_885_inst
    process(shl156_874, conv159_881) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl156_874, conv159_881, tmp_var);
      add160_886 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_903_inst
    process(shl162_892, conv165_899) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl162_892, conv165_899, tmp_var);
      add166_904 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_921_inst
    process(shl168_910, conv171_917) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_910, conv171_917, tmp_var);
      add172_922 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_591_inst
    process(conv70_586) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv70_586, type_cast_590_wire_constant, tmp_var);
      shl_592 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_609_inst
    process(add_604) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_604, type_cast_608_wire_constant, tmp_var);
      shl76_610 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_627_inst
    process(add80_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add80_622, type_cast_626_wire_constant, tmp_var);
      shl82_628 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_645_inst
    process(add86_640) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add86_640, type_cast_644_wire_constant, tmp_var);
      shl88_646 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_663_inst
    process(add92_658) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add92_658, type_cast_662_wire_constant, tmp_var);
      shl94_664 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_681_inst
    process(add98_676) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add98_676, type_cast_680_wire_constant, tmp_var);
      shl100_682 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_699_inst
    process(add104_694) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add104_694, type_cast_698_wire_constant, tmp_var);
      shl106_700 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_801_inst
    process(conv130_796) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv130_796, type_cast_800_wire_constant, tmp_var);
      shl132_802 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_819_inst
    process(add136_814) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add136_814, type_cast_818_wire_constant, tmp_var);
      shl138_820 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_837_inst
    process(add142_832) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add142_832, type_cast_836_wire_constant, tmp_var);
      shl144_838 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_855_inst
    process(add148_850) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add148_850, type_cast_854_wire_constant, tmp_var);
      shl150_856 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_873_inst
    process(add154_868) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add154_868, type_cast_872_wire_constant, tmp_var);
      shl156_874 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_891_inst
    process(add160_886) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add160_886, type_cast_890_wire_constant, tmp_var);
      shl162_892 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_909_inst
    process(add166_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_904, type_cast_908_wire_constant, tmp_var);
      shl168_910 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1016_inst
    process(tmp235_1011) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp235_1011, type_cast_1015_wire_constant, tmp_var);
      tmp236_1017 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_997_inst
    process(mul186_992) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul186_992, type_cast_996_wire_constant, tmp_var);
      cmp191204_998 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_554_inst
    process(tmp8_549) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp8_549, type_cast_553_wire_constant, tmp_var);
      tmp9_555 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_764_inst
    process(tmp16_759) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp16_759, type_cast_763_wire_constant, tmp_var);
      tmp17_765 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_129_inst
    process(inc_98, tmp1_125) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc_98, tmp1_125, tmp_var);
      cmp_130 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_239_inst
    process(inc22_201, tmp11_235) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc22_201, tmp11_235, tmp_var);
      cmp12_240 <= tmp_var; --
    end process;
    -- shared split operator group (69) : array_obj_ref_103_index_offset 
    ApIntAdd_group_69: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar268_102_scaled;
      array_obj_ref_103_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_103_index_offset_req_0;
      array_obj_ref_103_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_103_index_offset_req_1;
      array_obj_ref_103_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_69_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_69_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : array_obj_ref_1055_index_offset 
    ApIntAdd_group_70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1054_scaled;
      array_obj_ref_1055_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1055_index_offset_req_0;
      array_obj_ref_1055_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1055_index_offset_req_1;
      array_obj_ref_1055_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_70_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : array_obj_ref_206_index_offset 
    ApIntAdd_group_71: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar263_205_scaled;
      array_obj_ref_206_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_206_index_offset_req_0;
      array_obj_ref_206_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_206_index_offset_req_1;
      array_obj_ref_206_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_71_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_71_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_71",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : array_obj_ref_577_index_offset 
    ApIntAdd_group_72: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar250_576_scaled;
      array_obj_ref_577_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_577_index_offset_req_0;
      array_obj_ref_577_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_577_index_offset_req_1;
      array_obj_ref_577_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_72_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_72_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_72",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : array_obj_ref_787_index_offset 
    ApIntAdd_group_73: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar240_786_scaled;
      array_obj_ref_787_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_787_index_offset_req_0;
      array_obj_ref_787_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_787_index_offset_req_1;
      array_obj_ref_787_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_73_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_73_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_73",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100001",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared load operator group (0) : ptr_deref_407_load_0 ptr_deref_124_load_0 ptr_deref_383_load_0 ptr_deref_395_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_407_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_124_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_383_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_395_load_0_req_0;
      ptr_deref_407_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_124_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_383_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_395_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_407_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_124_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_383_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_395_load_0_req_1;
      ptr_deref_407_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_124_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_383_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_395_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_407_word_address_0 & ptr_deref_124_word_address_0 & ptr_deref_383_word_address_0 & ptr_deref_395_word_address_0;
      ptr_deref_407_data_0 <= data_out(127 downto 96);
      ptr_deref_124_data_0 <= data_out(95 downto 64);
      ptr_deref_383_data_0 <= data_out(63 downto 32);
      ptr_deref_395_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_433_load_0 ptr_deref_445_load_0 ptr_deref_457_load_0 ptr_deref_469_load_0 ptr_deref_234_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(34 downto 0);
      signal data_out: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= ptr_deref_433_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_445_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_457_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_469_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_234_load_0_req_0;
      ptr_deref_433_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_445_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_457_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_469_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_234_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= ptr_deref_433_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_445_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_457_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_469_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_234_load_0_req_1;
      ptr_deref_433_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_445_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_457_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_469_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_234_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_433_word_address_0 & ptr_deref_445_word_address_0 & ptr_deref_457_word_address_0 & ptr_deref_469_word_address_0 & ptr_deref_234_word_address_0;
      ptr_deref_433_data_0 <= data_out(159 downto 128);
      ptr_deref_445_data_0 <= data_out(127 downto 96);
      ptr_deref_457_data_0 <= data_out(95 downto 64);
      ptr_deref_469_data_0 <= data_out(63 downto 32);
      ptr_deref_234_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_981_load_0 ptr_deref_969_load_0 ptr_deref_957_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_981_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_969_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_957_load_0_req_0;
      ptr_deref_981_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_969_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_957_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_981_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_969_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_957_load_0_req_1;
      ptr_deref_981_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_969_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_957_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_981_word_address_0 & ptr_deref_969_word_address_0 & ptr_deref_957_word_address_0;
      ptr_deref_981_data_0 <= data_out(95 downto 64);
      ptr_deref_969_data_0 <= data_out(63 downto 32);
      ptr_deref_957_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : STORE_padding_313_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_padding_313_store_0_req_0;
      STORE_padding_313_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_padding_313_store_0_req_1;
      STORE_padding_313_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_padding_313_word_address_0;
      data_in <= STORE_padding_313_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1059_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1059_store_0_req_0;
      ptr_deref_1059_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1059_store_0_req_1;
      ptr_deref_1059_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1059_word_address_0;
      data_in <= ptr_deref_1059_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_49_store_0 ptr_deref_107_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_49_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_107_store_0_req_0;
      ptr_deref_49_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_107_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_49_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_107_store_0_req_1;
      ptr_deref_49_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_107_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_49_word_address_0 & ptr_deref_107_word_address_0;
      data_in <= ptr_deref_49_data_0 & ptr_deref_107_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_166_store_0 ptr_deref_217_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_166_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_217_store_0_req_0;
      ptr_deref_166_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_217_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_166_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_217_store_0_req_1;
      ptr_deref_166_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_217_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup3_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_166_word_address_0 & ptr_deref_217_word_address_0;
      data_in <= ptr_deref_166_data_0 & ptr_deref_217_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_279_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_279_store_0_req_0;
      ptr_deref_279_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_279_store_0_req_1;
      ptr_deref_279_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_279_word_address_0;
      data_in <= ptr_deref_279_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(15 downto 0),
          mtag => memory_space_8_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_332_store_0 ptr_deref_351_store_0 ptr_deref_370_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_332_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_351_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_370_store_0_req_0;
      ptr_deref_332_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_351_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_370_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_332_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_351_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_370_store_0_req_1;
      ptr_deref_332_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_351_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_370_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup5_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_332_word_address_0 & ptr_deref_351_word_address_0 & ptr_deref_370_word_address_0;
      data_in <= ptr_deref_332_data_0 & ptr_deref_351_data_0 & ptr_deref_370_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(6 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_714_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_714_store_0_req_0;
      ptr_deref_714_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_714_store_0_req_1;
      ptr_deref_714_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_714_word_address_0;
      data_in <= ptr_deref_714_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(13 downto 0),
          mdata => memory_space_4_sr_data(63 downto 0),
          mtag => memory_space_4_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_924_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_924_store_0_req_0;
      ptr_deref_924_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_924_store_0_req_1;
      ptr_deref_924_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup7_gI: SplitGuardInterface generic map(name => "StoreGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_924_word_address_0;
      data_in <= ptr_deref_924_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup7 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(10 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup7 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_612_inst RPIPE_ConvTranspose_input_pipe_666_inst RPIPE_ConvTranspose_input_pipe_648_inst RPIPE_ConvTranspose_input_pipe_630_inst RPIPE_ConvTranspose_input_pipe_894_inst RPIPE_ConvTranspose_input_pipe_684_inst RPIPE_ConvTranspose_input_pipe_840_inst RPIPE_ConvTranspose_input_pipe_702_inst RPIPE_ConvTranspose_input_pipe_791_inst RPIPE_ConvTranspose_input_pipe_912_inst RPIPE_ConvTranspose_input_pipe_581_inst RPIPE_ConvTranspose_input_pipe_858_inst RPIPE_ConvTranspose_input_pipe_876_inst RPIPE_ConvTranspose_input_pipe_594_inst RPIPE_ConvTranspose_input_pipe_804_inst RPIPE_ConvTranspose_input_pipe_822_inst RPIPE_ConvTranspose_input_pipe_36_inst RPIPE_ConvTranspose_input_pipe_60_inst RPIPE_ConvTranspose_input_pipe_132_inst RPIPE_ConvTranspose_input_pipe_210_inst RPIPE_ConvTranspose_input_pipe_251_inst RPIPE_ConvTranspose_input_pipe_283_inst RPIPE_ConvTranspose_input_pipe_317_inst RPIPE_ConvTranspose_input_pipe_336_inst RPIPE_ConvTranspose_input_pipe_355_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(199 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 24 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 24 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 24 downto 0);
      signal guard_vector : std_logic_vector( 24 downto 0);
      constant outBUFs : IntegerArray(24 downto 0) := (24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(24 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false);
      constant guardBuffering: IntegerArray(24 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2);
      -- 
    begin -- 
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_612_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_666_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_648_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_630_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_894_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_684_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_840_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_702_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_791_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_912_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_581_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_858_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_876_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_594_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_804_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_822_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_36_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_132_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_210_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_251_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_283_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_317_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_336_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_355_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_612_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_666_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_648_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_630_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_894_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_684_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_840_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_702_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_791_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_912_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_581_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_858_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_876_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_594_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_804_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_822_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_36_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_132_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_210_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_251_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_283_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_317_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_336_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_355_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_612_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_666_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_648_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_630_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_894_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_684_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_840_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_702_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_791_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_912_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_581_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_858_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_876_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_594_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_804_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_822_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_36_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_132_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_210_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_251_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_283_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_317_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_336_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_355_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_612_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_666_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_648_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_630_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_894_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_684_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_840_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_702_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_791_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_912_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_581_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_858_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_876_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_594_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_804_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_822_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_36_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_132_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_210_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_251_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_283_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_317_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_336_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_355_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      call77_613 <= data_out(199 downto 192);
      call95_667 <= data_out(191 downto 184);
      call89_649 <= data_out(183 downto 176);
      call83_631 <= data_out(175 downto 168);
      call163_895 <= data_out(167 downto 160);
      call101_685 <= data_out(159 downto 152);
      call145_841 <= data_out(151 downto 144);
      call107_703 <= data_out(143 downto 136);
      call129_792 <= data_out(135 downto 128);
      call169_913 <= data_out(127 downto 120);
      call69_582 <= data_out(119 downto 112);
      call151_859 <= data_out(111 downto 104);
      call157_877 <= data_out(103 downto 96);
      call72_595 <= data_out(95 downto 88);
      call133_805 <= data_out(87 downto 80);
      call139_823 <= data_out(79 downto 72);
      call_37 <= data_out(71 downto 64);
      call3228_61 <= data_out(63 downto 56);
      call3_133 <= data_out(55 downto 48);
      call15_211 <= data_out(47 downto 40);
      call29217_252 <= data_out(39 downto 32);
      call29_284 <= data_out(31 downto 24);
      call40_318 <= data_out(23 downto 16);
      call42_337 <= data_out(15 downto 8);
      call44_356 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 25, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 25,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_3266_start: Boolean;
  signal timer_CP_3266_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_1094_load_0_req_1 : boolean;
  signal LOAD_count_1094_load_0_ack_1 : boolean;
  signal LOAD_count_1094_load_0_req_0 : boolean;
  signal LOAD_count_1094_load_0_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_3266_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_3266_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_3266_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_3266_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_3266: Block -- control-path 
    signal timer_CP_3266_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_3266_elements(0) <= timer_CP_3266_start;
    timer_CP_3266_symbol <= timer_CP_3266_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_update_start_
      -- CP-element group 0: 	 assign_stmt_1095/LOAD_count_1094_sample_start_
      -- CP-element group 0: 	 assign_stmt_1095/$entry
      -- CP-element group 0: 	 $entry
      -- 
    cr_3298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_3266_elements(0), ack => LOAD_count_1094_load_0_req_1); -- 
    rr_3287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_3266_elements(0), ack => LOAD_count_1094_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_1095/LOAD_count_1094_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_1095/LOAD_count_1094_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_1095/LOAD_count_1094_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_1095/LOAD_count_1094_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1095/LOAD_count_1094_sample_completed_
      -- 
    ra_3288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_1094_load_0_ack_0, ack => timer_CP_3266_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_Update/LOAD_count_1094_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_Update/LOAD_count_1094_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_Update/LOAD_count_1094_Merge/merge_ack
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_Update/LOAD_count_1094_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_1095/LOAD_count_1094_update_completed_
      -- CP-element group 2: 	 assign_stmt_1095/$exit
      -- CP-element group 2: 	 $exit
      -- 
    ca_3299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_1094_load_0_ack_1, ack => timer_CP_3266_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_1094_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_1094_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_1094_word_address_0 <= "0";
    -- equivalence LOAD_count_1094_gather_scatter
    process(LOAD_count_1094_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_1094_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_1094_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_1094_load_0_req_0;
      LOAD_count_1094_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_1094_load_0_req_1;
      LOAD_count_1094_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_1094_word_address_0;
      LOAD_count_1094_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(5 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(5 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(41 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(119 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(5 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(5 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(191 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(11 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 21),
      memory_space_1_lr_tag => memory_space_1_lr_tag(83 downto 63),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 96),
      memory_space_1_lc_tag => memory_space_1_lc_tag(11 downto 9),
      memory_space_2_lr_req => memory_space_2_lr_req(3 downto 3),
      memory_space_2_lr_ack => memory_space_2_lr_ack(3 downto 3),
      memory_space_2_lr_addr => memory_space_2_lr_addr(27 downto 21),
      memory_space_2_lr_tag => memory_space_2_lr_tag(83 downto 63),
      memory_space_2_lc_req => memory_space_2_lc_req(3 downto 3),
      memory_space_2_lc_ack => memory_space_2_lc_ack(3 downto 3),
      memory_space_2_lc_data => memory_space_2_lc_data(127 downto 96),
      memory_space_2_lc_tag => memory_space_2_lc_tag(11 downto 9),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 21),
      memory_space_3_lr_tag => memory_space_3_lr_tag(79 downto 60),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(127 downto 96),
      memory_space_3_lc_tag => memory_space_3_lc_tag(7 downto 6),
      memory_space_4_lr_req => memory_space_4_lr_req(3 downto 3),
      memory_space_4_lr_ack => memory_space_4_lr_ack(3 downto 3),
      memory_space_4_lr_addr => memory_space_4_lr_addr(55 downto 42),
      memory_space_4_lr_tag => memory_space_4_lr_tag(75 downto 57),
      memory_space_4_lc_req => memory_space_4_lc_req(3 downto 3),
      memory_space_4_lc_ack => memory_space_4_lc_ack(3 downto 3),
      memory_space_4_lc_data => memory_space_4_lc_data(255 downto 192),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 3),
      memory_space_7_lr_req => memory_space_7_lr_req(3 downto 3),
      memory_space_7_lr_ack => memory_space_7_lr_ack(3 downto 3),
      memory_space_7_lr_addr => memory_space_7_lr_addr(3 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(75 downto 57),
      memory_space_7_lc_req => memory_space_7_lc_req(3 downto 3),
      memory_space_7_lc_ack => memory_space_7_lc_ack(3 downto 3),
      memory_space_7_lc_data => memory_space_7_lc_data(63 downto 48),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 3),
      memory_space_8_lr_req => memory_space_8_lr_req(3 downto 3),
      memory_space_8_lr_ack => memory_space_8_lr_ack(3 downto 3),
      memory_space_8_lr_addr => memory_space_8_lr_addr(3 downto 3),
      memory_space_8_lr_tag => memory_space_8_lr_tag(79 downto 60),
      memory_space_8_lc_req => memory_space_8_lc_req(3 downto 3),
      memory_space_8_lc_ack => memory_space_8_lc_ack(3 downto 3),
      memory_space_8_lc_data => memory_space_8_lc_data(63 downto 48),
      memory_space_8_lc_tag => memory_space_8_lc_tag(7 downto 6),
      memory_space_6_sr_req => memory_space_6_sr_req(3 downto 3),
      memory_space_6_sr_ack => memory_space_6_sr_ack(3 downto 3),
      memory_space_6_sr_addr => memory_space_6_sr_addr(55 downto 42),
      memory_space_6_sr_data => memory_space_6_sr_data(255 downto 192),
      memory_space_6_sr_tag => memory_space_6_sr_tag(75 downto 57),
      memory_space_6_sc_req => memory_space_6_sc_req(3 downto 3),
      memory_space_6_sc_ack => memory_space_6_sc_ack(3 downto 3),
      memory_space_6_sc_tag => memory_space_6_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(20 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(62 downto 42),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(95 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(8 downto 6),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(20 downto 14),
      memory_space_2_lr_tag => memory_space_2_lr_tag(62 downto 42),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(95 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(8 downto 6),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(20 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(59 downto 40),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(95 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(5 downto 4),
      memory_space_4_lr_req => memory_space_4_lr_req(2 downto 2),
      memory_space_4_lr_ack => memory_space_4_lr_ack(2 downto 2),
      memory_space_4_lr_addr => memory_space_4_lr_addr(41 downto 28),
      memory_space_4_lr_tag => memory_space_4_lr_tag(56 downto 38),
      memory_space_4_lc_req => memory_space_4_lc_req(2 downto 2),
      memory_space_4_lc_ack => memory_space_4_lc_ack(2 downto 2),
      memory_space_4_lc_data => memory_space_4_lc_data(191 downto 128),
      memory_space_4_lc_tag => memory_space_4_lc_tag(2 downto 2),
      memory_space_7_lr_req => memory_space_7_lr_req(2 downto 2),
      memory_space_7_lr_ack => memory_space_7_lr_ack(2 downto 2),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 2),
      memory_space_7_lr_tag => memory_space_7_lr_tag(56 downto 38),
      memory_space_7_lc_req => memory_space_7_lc_req(2 downto 2),
      memory_space_7_lc_ack => memory_space_7_lc_ack(2 downto 2),
      memory_space_7_lc_data => memory_space_7_lc_data(47 downto 32),
      memory_space_7_lc_tag => memory_space_7_lc_tag(2 downto 2),
      memory_space_8_lr_req => memory_space_8_lr_req(2 downto 2),
      memory_space_8_lr_ack => memory_space_8_lr_ack(2 downto 2),
      memory_space_8_lr_addr => memory_space_8_lr_addr(2 downto 2),
      memory_space_8_lr_tag => memory_space_8_lr_tag(59 downto 40),
      memory_space_8_lc_req => memory_space_8_lc_req(2 downto 2),
      memory_space_8_lc_ack => memory_space_8_lc_ack(2 downto 2),
      memory_space_8_lc_data => memory_space_8_lc_data(47 downto 32),
      memory_space_8_lc_tag => memory_space_8_lc_tag(5 downto 4),
      memory_space_6_sr_req => memory_space_6_sr_req(2 downto 2),
      memory_space_6_sr_ack => memory_space_6_sr_ack(2 downto 2),
      memory_space_6_sr_addr => memory_space_6_sr_addr(41 downto 28),
      memory_space_6_sr_data => memory_space_6_sr_data(191 downto 128),
      memory_space_6_sr_tag => memory_space_6_sr_tag(56 downto 38),
      memory_space_6_sc_req => memory_space_6_sc_req(2 downto 2),
      memory_space_6_sc_ack => memory_space_6_sc_ack(2 downto 2),
      memory_space_6_sc_tag => memory_space_6_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 7),
      memory_space_1_lr_tag => memory_space_1_lr_tag(41 downto 21),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 3),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 7),
      memory_space_2_lr_tag => memory_space_2_lr_tag(41 downto 21),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 3),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 7),
      memory_space_3_lr_tag => memory_space_3_lr_tag(39 downto 20),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 32),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 2),
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(27 downto 14),
      memory_space_4_lr_tag => memory_space_4_lr_tag(37 downto 19),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(127 downto 64),
      memory_space_4_lc_tag => memory_space_4_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(37 downto 19),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 16),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 1),
      memory_space_8_lr_req => memory_space_8_lr_req(1 downto 1),
      memory_space_8_lr_ack => memory_space_8_lr_ack(1 downto 1),
      memory_space_8_lr_addr => memory_space_8_lr_addr(1 downto 1),
      memory_space_8_lr_tag => memory_space_8_lr_tag(39 downto 20),
      memory_space_8_lc_req => memory_space_8_lc_req(1 downto 1),
      memory_space_8_lc_ack => memory_space_8_lc_ack(1 downto 1),
      memory_space_8_lc_data => memory_space_8_lc_data(31 downto 16),
      memory_space_8_lc_tag => memory_space_8_lc_tag(3 downto 2),
      memory_space_6_sr_req => memory_space_6_sr_req(1 downto 1),
      memory_space_6_sr_ack => memory_space_6_sr_ack(1 downto 1),
      memory_space_6_sr_addr => memory_space_6_sr_addr(27 downto 14),
      memory_space_6_sr_data => memory_space_6_sr_data(127 downto 64),
      memory_space_6_sr_tag => memory_space_6_sr_tag(37 downto 19),
      memory_space_6_sc_req => memory_space_6_sc_req(1 downto 1),
      memory_space_6_sc_ack => memory_space_6_sc_ack(1 downto 1),
      memory_space_6_sc_tag => memory_space_6_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(20 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(2 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(6 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(19 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(13 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(18 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(63 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(18 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(0 downto 0),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(0 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(19 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(15 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(1 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(13 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(63 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(4 downto 4),
      memory_space_3_lr_ack => memory_space_3_lr_ack(4 downto 4),
      memory_space_3_lr_addr => memory_space_3_lr_addr(34 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(99 downto 80),
      memory_space_3_lc_req => memory_space_3_lc_req(4 downto 4),
      memory_space_3_lc_ack => memory_space_3_lc_ack(4 downto 4),
      memory_space_3_lc_data => memory_space_3_lc_data(159 downto 128),
      memory_space_3_lc_tag => memory_space_3_lc_tag(9 downto 8),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(13 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(34 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(104 downto 84),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(159 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(14 downto 12),
      memory_space_2_lr_req => memory_space_2_lr_req(4 downto 4),
      memory_space_2_lr_ack => memory_space_2_lr_ack(4 downto 4),
      memory_space_2_lr_addr => memory_space_2_lr_addr(34 downto 28),
      memory_space_2_lr_tag => memory_space_2_lr_tag(104 downto 84),
      memory_space_2_lc_req => memory_space_2_lc_req(4 downto 4),
      memory_space_2_lc_ack => memory_space_2_lc_ack(4 downto 4),
      memory_space_2_lc_data => memory_space_2_lc_data(159 downto 128),
      memory_space_2_lc_tag => memory_space_2_lc_tag(14 downto 12),
      memory_space_3_lr_req => memory_space_3_lr_req(5 downto 5),
      memory_space_3_lr_ack => memory_space_3_lr_ack(5 downto 5),
      memory_space_3_lr_addr => memory_space_3_lr_addr(41 downto 35),
      memory_space_3_lr_tag => memory_space_3_lr_tag(119 downto 100),
      memory_space_3_lc_req => memory_space_3_lc_req(5 downto 5),
      memory_space_3_lc_ack => memory_space_3_lc_ack(5 downto 5),
      memory_space_3_lc_data => memory_space_3_lc_data(191 downto 160),
      memory_space_3_lc_tag => memory_space_3_lc_tag(11 downto 10),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(20 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(6 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(19 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(13 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(63 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(18 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(10 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(0 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(4 downto 4),
      memory_space_6_sr_ack => memory_space_6_sr_ack(4 downto 4),
      memory_space_6_sr_addr => memory_space_6_sr_addr(69 downto 56),
      memory_space_6_sr_data => memory_space_6_sr_data(319 downto 256),
      memory_space_6_sr_tag => memory_space_6_sr_tag(94 downto 76),
      memory_space_6_sc_req => memory_space_6_sc_req(4 downto 4),
      memory_space_6_sc_ack => memory_space_6_sc_ack(4 downto 4),
      memory_space_6_sc_tag => memory_space_6_sc_tag(4 downto 4),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(18 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(0 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(15 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(19 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 6,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_5: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
