-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    num_cont : in  std_logic_vector(15 downto 0);
    row1 : in  std_logic_vector(15 downto 0);
    col1 : in  std_logic_vector(15 downto 0);
    rk1 : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal num_cont_buffer :  std_logic_vector(15 downto 0);
  signal num_cont_update_enable: Boolean;
  signal row1_buffer :  std_logic_vector(15 downto 0);
  signal row1_update_enable: Boolean;
  signal col1_buffer :  std_logic_vector(15 downto 0);
  signal col1_update_enable: Boolean;
  signal rk1_buffer :  std_logic_vector(15 downto 0);
  signal rk1_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_44_branch_req_0 : boolean;
  signal phi_stmt_46_ack_0 : boolean;
  signal phi_stmt_46_req_1 : boolean;
  signal phi_stmt_46_req_0 : boolean;
  signal n_address_280_50_buf_req_0 : boolean;
  signal n_address_280_50_buf_ack_0 : boolean;
  signal n_address_280_50_buf_req_1 : boolean;
  signal n_address_280_50_buf_ack_1 : boolean;
  signal phi_stmt_51_req_1 : boolean;
  signal phi_stmt_51_req_0 : boolean;
  signal phi_stmt_51_ack_0 : boolean;
  signal n_word_start_269_56_buf_req_0 : boolean;
  signal n_word_start_269_56_buf_ack_0 : boolean;
  signal n_word_start_269_56_buf_req_1 : boolean;
  signal n_word_start_269_56_buf_ack_1 : boolean;
  signal n_winr_209_68_buf_req_1 : boolean;
  signal n_winr_209_68_buf_ack_1 : boolean;
  signal phi_stmt_57_req_1 : boolean;
  signal phi_stmt_57_req_0 : boolean;
  signal phi_stmt_57_ack_0 : boolean;
  signal nl_start_35_59_buf_req_0 : boolean;
  signal nl_start_35_59_buf_ack_0 : boolean;
  signal nl_start_35_59_buf_req_1 : boolean;
  signal nl_start_35_59_buf_ack_1 : boolean;
  signal n_left_288_60_buf_req_0 : boolean;
  signal n_left_288_60_buf_ack_0 : boolean;
  signal n_left_288_60_buf_req_1 : boolean;
  signal n_left_288_60_buf_ack_1 : boolean;
  signal phi_stmt_61_req_1 : boolean;
  signal phi_stmt_61_req_0 : boolean;
  signal phi_stmt_61_ack_0 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal n_blk_308_65_buf_req_0 : boolean;
  signal n_blk_308_65_buf_ack_0 : boolean;
  signal n_blk_308_65_buf_req_1 : boolean;
  signal n_blk_308_65_buf_ack_1 : boolean;
  signal phi_stmt_66_req_0 : boolean;
  signal phi_stmt_66_req_1 : boolean;
  signal phi_stmt_66_ack_0 : boolean;
  signal n_winr_209_68_buf_req_0 : boolean;
  signal n_winr_209_68_buf_ack_0 : boolean;
  signal WPIPE_input_pipe1_167_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_167_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_167_inst_ack_1 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_req_0 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_ack_0 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_req_1 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_ack_1 : boolean;
  signal phi_stmt_71_req_0 : boolean;
  signal phi_stmt_71_req_1 : boolean;
  signal phi_stmt_71_ack_0 : boolean;
  signal n_col_222_73_buf_req_0 : boolean;
  signal n_col_222_73_buf_ack_0 : boolean;
  signal n_col_222_73_buf_req_1 : boolean;
  signal n_col_222_73_buf_ack_1 : boolean;
  signal phi_stmt_76_req_0 : boolean;
  signal phi_stmt_76_req_1 : boolean;
  signal phi_stmt_76_ack_0 : boolean;
  signal n_row_234_78_buf_req_0 : boolean;
  signal n_row_234_78_buf_ack_0 : boolean;
  signal n_row_234_78_buf_req_1 : boolean;
  signal n_row_234_78_buf_ack_1 : boolean;
  signal array_obj_ref_133_index_offset_req_0 : boolean;
  signal array_obj_ref_133_index_offset_ack_0 : boolean;
  signal array_obj_ref_133_index_offset_req_1 : boolean;
  signal array_obj_ref_133_index_offset_ack_1 : boolean;
  signal addr_of_134_final_reg_req_0 : boolean;
  signal addr_of_134_final_reg_ack_0 : boolean;
  signal addr_of_134_final_reg_req_1 : boolean;
  signal addr_of_134_final_reg_ack_1 : boolean;
  signal ptr_deref_138_load_0_req_0 : boolean;
  signal ptr_deref_138_load_0_ack_0 : boolean;
  signal ptr_deref_138_load_0_req_1 : boolean;
  signal ptr_deref_138_load_0_ack_1 : boolean;
  signal slice_142_inst_req_0 : boolean;
  signal slice_142_inst_ack_0 : boolean;
  signal slice_142_inst_req_1 : boolean;
  signal slice_142_inst_ack_1 : boolean;
  signal slice_146_inst_req_0 : boolean;
  signal slice_146_inst_ack_0 : boolean;
  signal slice_146_inst_req_1 : boolean;
  signal slice_146_inst_ack_1 : boolean;
  signal slice_150_inst_req_0 : boolean;
  signal slice_150_inst_ack_0 : boolean;
  signal slice_150_inst_req_1 : boolean;
  signal slice_150_inst_ack_1 : boolean;
  signal slice_154_inst_req_0 : boolean;
  signal slice_154_inst_ack_0 : boolean;
  signal slice_154_inst_req_1 : boolean;
  signal slice_154_inst_ack_1 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_req_0 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_ack_0 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_req_1 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_160_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_160_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_160_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_160_inst_ack_1 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_req_0 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_ack_0 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_req_1 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_167_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_174_inst_ack_1 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_req_0 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_ack_0 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_req_1 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_181_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_181_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_181_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_181_inst_ack_1 : boolean;
  signal do_while_stmt_44_branch_ack_0 : boolean;
  signal do_while_stmt_44_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= num_cont;
  num_cont_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= row1;
  row1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= col1;
  col1_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= rk1;
  rk1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= ct;
  ct_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43__exit__
      -- CP-element group 0: 	 branch_block_stmt_26/do_while_stmt_44__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_26/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/branch_block_stmt_26__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	207 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_26/$exit
      -- CP-element group 1: 	 branch_block_stmt_26/branch_block_stmt_26__exit__
      -- CP-element group 1: 	 branch_block_stmt_26/do_while_stmt_44__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(207);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_26/do_while_stmt_44/$entry
      -- CP-element group 2: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	207 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_26/do_while_stmt_44/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	205 
    -- CP-element group 5: 	206 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/condition_done
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	204 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_26/do_while_stmt_44/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(204);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	77 
    -- CP-element group 7: 	135 
    -- CP-element group 7: 	116 
    -- CP-element group 7: 	58 
    -- CP-element group 7: 	98 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	100 
    -- CP-element group 8: 	137 
    -- CP-element group 8: 	118 
    -- CP-element group 8: 	79 
    -- CP-element group 8: 	60 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	203 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	111 
    -- CP-element group 9: 	92 
    -- CP-element group 9: 	72 
    -- CP-element group 9: 	112 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	149 
    -- CP-element group 9: 	130 
    -- CP-element group 9: 	54 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	93 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	203 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_44_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(203) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	71 
    -- CP-element group 11: 	111 
    -- CP-element group 11: 	92 
    -- CP-element group 11: 	129 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	73 
    -- CP-element group 11: 	94 
    -- CP-element group 11: 	131 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= access_T_CP_0_elements(71) & access_T_CP_0_elements(111) & access_T_CP_0_elements(92) & access_T_CP_0_elements(129) & access_T_CP_0_elements(53) & access_T_CP_0_elements(15) & access_T_CP_0_elements(34) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	113 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	95 
    -- CP-element group 12: 	74 
    -- CP-element group 12: 	132 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	204 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	71 
    -- CP-element group 12: 	111 
    -- CP-element group 12: 	92 
    -- CP-element group 12: 	129 
    -- CP-element group 12: 	53 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(113) & access_T_CP_0_elements(56) & access_T_CP_0_elements(95) & access_T_CP_0_elements(74) & access_T_CP_0_elements(132) & access_T_CP_0_elements(18) & access_T_CP_0_elements(37);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	72 
    -- CP-element group 13: 	112 
    -- CP-element group 13: 	130 
    -- CP-element group 13: 	54 
    -- CP-element group 13: 	93 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	75 
    -- CP-element group 13: 	96 
    -- CP-element group 13: 	114 
    -- CP-element group 13: 	133 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(72) & access_T_CP_0_elements(112) & access_T_CP_0_elements(130) & access_T_CP_0_elements(54) & access_T_CP_0_elements(93) & access_T_CP_0_elements(16) & access_T_CP_0_elements(35);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	97 
    -- CP-element group 14: 	76 
    -- CP-element group 14: 	115 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	134 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(97) & access_T_CP_0_elements(76) & access_T_CP_0_elements(115) & access_T_CP_0_elements(57) & access_T_CP_0_elements(134) & access_T_CP_0_elements(20) & access_T_CP_0_elements(39);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	151 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start__ps
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start__ps
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(13);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	151 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (15) 
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resized_1
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scaled_1
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_computed_1
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/index_resize_req
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/index_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/scale_rename_req
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/scale_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/req
      -- 
    req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => array_obj_ref_133_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req_ps
      -- 
    phi_stmt_46_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_46_req_1); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_trigger
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req_ps
      -- 
    phi_stmt_46_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => phi_stmt_46_req_0); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack_ps
      -- 
    phi_stmt_46_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_46_ack_0, ack => access_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_start_
      -- 
    -- Element group access_T_CP_0_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_completed__ps
      -- 
    access_T_CP_0_elements(28) <= access_T_CP_0_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(27), ack => access_T_CP_0_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/req
      -- 
    req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(30), ack => n_address_280_50_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_start_
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/req
      -- 
    req_76_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_76_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(31), ack => n_address_280_50_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/ack
      -- 
    ack_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_280_50_buf_ack_0, ack => access_T_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/ack
      -- 
    ack_77_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_280_50_buf_ack_1, ack => access_T_CP_0_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_start_
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	198 
    -- CP-element group 35: 	191 
    -- CP-element group 35: 	177 
    -- CP-element group 35: 	184 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_start_
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(198) & access_T_CP_0_elements(191) & access_T_CP_0_elements(177) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: 	196 
    -- CP-element group 39: 	189 
    -- CP-element group 39: 	175 
    -- CP-element group 39: 	182 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_sample_req_ps
      -- 
    phi_stmt_51_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_51_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_51_req_1); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_sample_req_ps
      -- 
    phi_stmt_51_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_51_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_51_req_0); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_phi_mux_ack_ps
      -- 
    phi_stmt_51_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_51_ack_0, ack => access_T_CP_0_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_start_
      -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_completed__ps
      -- 
    access_T_CP_0_elements(47) <= access_T_CP_0_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(46), ack => access_T_CP_0_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/req
      -- 
    req_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(49), ack => n_word_start_269_56_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_start_
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/req
      -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(50), ack => n_word_start_269_56_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/ack
      -- 
    ack_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_269_56_buf_ack_0, ack => access_T_CP_0_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_269_56_buf_ack_1, ack => access_T_CP_0_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	11 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_start_
      -- 
    access_T_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_start_
      -- 
    access_T_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(57);
      gj_access_T_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_start__ps
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(11);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	14 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	54 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(57) is bound as output of CP function.
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	7 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_trigger
      -- 
    access_T_CP_0_elements(58) <= access_T_CP_0_elements(7);
    -- CP-element group 59:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_sample_req
      -- CP-element group 59: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_sample_req_ps
      -- 
    phi_stmt_57_loopback_sample_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_loopback_sample_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(59), ack => phi_stmt_57_req_1); -- 
    -- Element group access_T_CP_0_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	8 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_trigger
      -- 
    access_T_CP_0_elements(60) <= access_T_CP_0_elements(8);
    -- CP-element group 61:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_sample_req
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_sample_req_ps
      -- 
    phi_stmt_57_entry_sample_req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_entry_sample_req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(61), ack => phi_stmt_57_req_0); -- 
    -- Element group access_T_CP_0_elements(61) is bound as output of CP function.
    -- CP-element group 62:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_phi_mux_ack
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_phi_mux_ack_ps
      -- 
    phi_stmt_57_phi_mux_ack_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_57_ack_0, ack => access_T_CP_0_elements(62)); -- 
    -- CP-element group 63:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_start__ps
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/req
      -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(63), ack => nl_start_35_59_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_start__ps
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_start_
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/req
      -- 
    req_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => nl_start_35_59_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_completed__ps
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_35_59_buf_ack_0, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/ack
      -- 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_35_59_buf_ack_1, ack => access_T_CP_0_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/req
      -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(67), ack => n_left_288_60_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_start__ps
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_start_
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(68), ack => n_left_288_60_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/ack
      -- 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_288_60_buf_ack_0, ack => access_T_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/ack
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_288_60_buf_ack_1, ack => access_T_CP_0_elements(70)); -- 
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	12 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	11 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_start_
      -- 
    access_T_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	9 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	198 
    -- CP-element group 72: 	191 
    -- CP-element group 72: 	184 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	13 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_start_
      -- 
    access_T_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(198) & access_T_CP_0_elements(191) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	11 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_start__ps
      -- 
    access_T_CP_0_elements(73) <= access_T_CP_0_elements(11);
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	12 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(74) is bound as output of CP function.
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	13 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_start__ps
      -- 
    access_T_CP_0_elements(75) <= access_T_CP_0_elements(13);
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	14 
    -- CP-element group 76: 	196 
    -- CP-element group 76: 	189 
    -- CP-element group 76: 	182 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(76) is bound as output of CP function.
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	7 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_trigger
      -- 
    access_T_CP_0_elements(77) <= access_T_CP_0_elements(7);
    -- CP-element group 78:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_sample_req
      -- CP-element group 78: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_sample_req_ps
      -- 
    phi_stmt_61_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_61_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(78), ack => phi_stmt_61_req_1); -- 
    -- Element group access_T_CP_0_elements(78) is bound as output of CP function.
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	8 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_trigger
      -- 
    access_T_CP_0_elements(79) <= access_T_CP_0_elements(8);
    -- CP-element group 80:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_sample_req
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_sample_req_ps
      -- 
    phi_stmt_61_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_61_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(80), ack => phi_stmt_61_req_0); -- 
    -- Element group access_T_CP_0_elements(80) is bound as output of CP function.
    -- CP-element group 81:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_phi_mux_ack
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_phi_mux_ack_ps
      -- 
    phi_stmt_61_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_61_ack_0, ack => access_T_CP_0_elements(81)); -- 
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/rr
      -- 
    rr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(84), ack => type_cast_64_inst_req_0); -- 
    access_T_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(82) & access_T_CP_0_elements(86);
      gj_access_T_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_start_
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/cr
      -- 
    cr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(85), ack => type_cast_64_inst_req_1); -- 
    access_T_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(83) & access_T_CP_0_elements(87);
      gj_access_T_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/ra
      -- 
    ra_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/ca
      -- 
    ca_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => access_T_CP_0_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_start__ps
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/req
      -- 
    req_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(88), ack => n_blk_308_65_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_start__ps
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_start_
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/req
      -- 
    req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(89), ack => n_blk_308_65_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/ack
      -- 
    ack_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_308_65_buf_ack_0, ack => access_T_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/ack
      -- 
    ack_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_308_65_buf_ack_1, ack => access_T_CP_0_elements(91)); -- 
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	9 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	12 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	11 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_start_
      -- 
    access_T_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	9 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	97 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	13 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_start_
      -- 
    access_T_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(97);
      gj_access_T_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	11 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_start__ps
      -- 
    access_T_CP_0_elements(94) <= access_T_CP_0_elements(11);
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	12 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(95) is bound as output of CP function.
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	13 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_start__ps
      -- 
    access_T_CP_0_elements(96) <= access_T_CP_0_elements(13);
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	14 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	93 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(97) is bound as output of CP function.
    -- CP-element group 98:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	7 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_trigger
      -- 
    access_T_CP_0_elements(98) <= access_T_CP_0_elements(7);
    -- CP-element group 99:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_sample_req
      -- CP-element group 99: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_sample_req_ps
      -- 
    phi_stmt_66_loopback_sample_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_loopback_sample_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(99), ack => phi_stmt_66_req_0); -- 
    -- Element group access_T_CP_0_elements(99) is bound as output of CP function.
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	8 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_trigger
      -- 
    access_T_CP_0_elements(100) <= access_T_CP_0_elements(8);
    -- CP-element group 101:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_sample_req
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_sample_req_ps
      -- 
    phi_stmt_66_entry_sample_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_entry_sample_req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(101), ack => phi_stmt_66_req_1); -- 
    -- Element group access_T_CP_0_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_phi_mux_ack
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_phi_mux_ack_ps
      -- 
    phi_stmt_66_phi_mux_ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_66_ack_0, ack => access_T_CP_0_elements(102)); -- 
    -- CP-element group 103:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_start__ps
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/req
      -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(103), ack => n_winr_209_68_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/req
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_start__ps
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_start_
      -- 
    req_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(104), ack => n_winr_209_68_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_completed__ps
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_209_68_buf_ack_0, ack => access_T_CP_0_elements(105)); -- 
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/ack
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_completed_
      -- 
    ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_209_68_buf_ack_1, ack => access_T_CP_0_elements(106)); -- 
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_start__ps
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_start__ps
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_start_
      -- 
    -- Element group access_T_CP_0_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_completed__ps
      -- 
    access_T_CP_0_elements(109) <= access_T_CP_0_elements(110);
    -- CP-element group 110:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	109 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(110) is a control-delay.
    cp_element_110_delay: control_delay_element  generic map(name => " 110_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(108), ack => access_T_CP_0_elements(110), clk => clk, reset =>reset);
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	9 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	12 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	11 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_start_
      -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	9 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	115 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	13 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_start_
      -- 
    access_T_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(115);
      gj_access_T_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	12 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	13 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_start__ps
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(13);
    -- CP-element group 115:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	14 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	112 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	7 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_trigger
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(7);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_sample_req
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_sample_req_ps
      -- 
    phi_stmt_71_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(117), ack => phi_stmt_71_req_0); -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	8 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_trigger
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(8);
    -- CP-element group 119:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_sample_req
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_sample_req_ps
      -- 
    phi_stmt_71_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => phi_stmt_71_req_1); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_phi_mux_ack
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_phi_mux_ack_ps
      -- 
    phi_stmt_71_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_71_ack_0, ack => access_T_CP_0_elements(120)); -- 
    -- CP-element group 121:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_sample_start__ps
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Sample/req
      -- 
    req_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(121), ack => n_col_222_73_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (4) 
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_update_start__ps
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_update_start_
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Update/req
      -- 
    req_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(122), ack => n_col_222_73_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_sample_completed__ps
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Sample/ack
      -- 
    ack_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_222_73_buf_ack_0, ack => access_T_CP_0_elements(123)); -- 
    -- CP-element group 124:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_update_completed__ps
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Update/ack
      -- 
    ack_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_222_73_buf_ack_1, ack => access_T_CP_0_elements(124)); -- 
    -- CP-element group 125:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_sample_completed__ps
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_update_start_
      -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_update_completed__ps
      -- 
    access_T_CP_0_elements(127) <= access_T_CP_0_elements(128);
    -- CP-element group 128:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	127 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(128) is a control-delay.
    cp_element_128_delay: control_delay_element  generic map(name => " 128_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(126), ack => access_T_CP_0_elements(128), clk => clk, reset =>reset);
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	12 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	11 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_start_
      -- 
    access_T_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	9 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	134 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	13 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_start_
      -- 
    access_T_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	11 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_start__ps
      -- 
    access_T_CP_0_elements(131) <= access_T_CP_0_elements(11);
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	12 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	13 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_start__ps
      -- 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(13);
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	14 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	130 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	7 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(7);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_sample_req
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_sample_req_ps
      -- 
    phi_stmt_76_loopback_sample_req_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_loopback_sample_req_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_76_req_0); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	8 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_trigger
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(8);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_sample_req
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_sample_req_ps
      -- 
    phi_stmt_76_entry_sample_req_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_entry_sample_req_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => phi_stmt_76_req_1); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_phi_mux_ack
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_phi_mux_ack_ps
      -- 
    phi_stmt_76_phi_mux_ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_76_ack_0, ack => access_T_CP_0_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Sample/req
      -- 
    req_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(140), ack => n_row_234_78_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_update_start_
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Update/req
      -- 
    req_352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(141), ack => n_row_234_78_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_sample_completed__ps
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Sample/ack
      -- 
    ack_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_234_78_buf_ack_0, ack => access_T_CP_0_elements(142)); -- 
    -- CP-element group 143:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_update_completed__ps
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Update/ack
      -- 
    ack_353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_234_78_buf_ack_1, ack => access_T_CP_0_elements(143)); -- 
    -- CP-element group 144:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_sample_start__ps
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_sample_completed__ps
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_update_start__ps
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_update_start_
      -- 
    -- Element group access_T_CP_0_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_update_completed__ps
      -- 
    access_T_CP_0_elements(146) <= access_T_CP_0_elements(147);
    -- CP-element group 147:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(147) is a control-delay.
    cp_element_147_delay: control_delay_element  generic map(name => " 147_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(145), ack => access_T_CP_0_elements(147), clk => clk, reset =>reset);
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	152 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/$entry
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/req
      -- 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => addr_of_134_final_reg_req_0); -- 
    access_T_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(152) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	9 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	157 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_update_start_
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/req
      -- 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(149), ack => addr_of_134_final_reg_req_1); -- 
    access_T_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_update_start
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/req
      -- 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => array_obj_ref_133_index_offset_req_1); -- 
    access_T_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	20 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	204 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	16 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_sample_complete
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/ack
      -- 
    ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_133_index_offset_ack_0, ack => access_T_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	148 
    -- CP-element group 152:  members (8) 
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_root_address_calculated
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_offset_calculated
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/$entry
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/sum_rename_req
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/sum_rename_ack
      -- 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_133_index_offset_ack_1, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/$exit
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/ack
      -- 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_134_final_reg_ack_0, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	149 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (19) 
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/root_register_ack
      -- 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_134_final_reg_ack_1, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/rr
      -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => ptr_deref_138_load_0_req_0); -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(154) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	169 
    -- CP-element group 156: 	173 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	165 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_update_start_
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/cr
      -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => ptr_deref_138_load_0_req_1); -- 
    access_T_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(169) & access_T_CP_0_elements(173) & access_T_CP_0_elements(161) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	149 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/ra
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_0, ack => access_T_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	167 
    -- CP-element group 158: 	171 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	163 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/ca
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/$entry
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/merge_req
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/merge_ack
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_1, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/rr
      -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(159), ack => slice_142_inst_req_0); -- 
    access_T_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(161);
      gj_access_T_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	180 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_update_start_
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/cr
      -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(160), ack => slice_142_inst_req_1); -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_0, ack => access_T_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	179 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/ca
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_1, ack => access_T_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/rr
      -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => slice_146_inst_req_0); -- 
    access_T_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	187 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_update_start_
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/cr
      -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(164), ack => slice_146_inst_req_1); -- 
    access_T_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	156 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/ra
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_0, ack => access_T_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	186 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/ca
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_1, ack => access_T_CP_0_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	158 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/rr
      -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => slice_150_inst_req_0); -- 
    access_T_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	194 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_update_start_
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/cr
      -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(168), ack => slice_150_inst_req_1); -- 
    access_T_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	156 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/ra
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_0, ack => access_T_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	193 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/ca
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_1, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	158 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/rr
      -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(171), ack => slice_154_inst_req_0); -- 
    access_T_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	201 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_update_start_
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/cr
      -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => slice_154_inst_req_1); -- 
    access_T_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	156 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/ra
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_0, ack => access_T_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	200 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/ca
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_1, ack => access_T_CP_0_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	39 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(175), ack => W_c1_156_delayed_14_0_156_inst_req_0); -- 
    access_T_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(39) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	180 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_update_start_
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/req
      -- 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => W_c1_156_delayed_14_0_156_inst_req_1); -- 
    access_T_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	35 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_156_delayed_14_0_156_inst_ack_0, ack => access_T_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/ack
      -- 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_156_delayed_14_0_156_inst_ack_1, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: 	162 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	202 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/req
      -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(179), ack => WPIPE_input_pipe1_160_inst_req_0); -- 
    access_T_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(178) & access_T_CP_0_elements(162) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	176 
    -- CP-element group 180: 	160 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_update_start_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/req
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_160_inst_ack_0, ack => access_T_CP_0_elements(180)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => WPIPE_input_pipe1_160_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_160_inst_ack_1, ack => access_T_CP_0_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	76 
    -- CP-element group 182: 	39 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/req
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => W_c2_160_delayed_14_0_163_inst_req_0); -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(76) & access_T_CP_0_elements(39) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	187 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_update_start_
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(183), ack => W_c2_160_delayed_14_0_163_inst_req_1); -- 
    access_T_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	72 
    -- CP-element group 184: 	35 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_160_delayed_14_0_163_inst_ack_0, ack => access_T_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_160_delayed_14_0_163_inst_ack_1, ack => access_T_CP_0_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: 	166 
    -- CP-element group 186: 	181 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/req
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(186), ack => WPIPE_input_pipe1_167_inst_req_0); -- 
    access_T_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(185) & access_T_CP_0_elements(166) & access_T_CP_0_elements(181) & access_T_CP_0_elements(188);
      gj_access_T_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	183 
    -- CP-element group 187: 	164 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/req
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_update_start_
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/$exit
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_167_inst_ack_0, ack => access_T_CP_0_elements(187)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(187), ack => WPIPE_input_pipe1_167_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_update_completed_
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_167_inst_ack_1, ack => access_T_CP_0_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	76 
    -- CP-element group 189: 	39 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => W_c3_164_delayed_14_0_170_inst_req_0); -- 
    access_T_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(76) & access_T_CP_0_elements(39) & access_T_CP_0_elements(191);
      gj_access_T_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_update_start_
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/req
      -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => W_c3_164_delayed_14_0_170_inst_req_1); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	72 
    -- CP-element group 191: 	35 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_164_delayed_14_0_170_inst_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/ack
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_164_delayed_14_0_170_inst_ack_1, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	192 
    -- CP-element group 193: 	170 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/req
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => WPIPE_input_pipe1_174_inst_req_0); -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(188) & access_T_CP_0_elements(192) & access_T_CP_0_elements(170) & access_T_CP_0_elements(195);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	168 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_update_start_
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/req
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_174_inst_ack_0, ack => access_T_CP_0_elements(194)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(194), ack => WPIPE_input_pipe1_174_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/ack
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_174_inst_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	76 
    -- CP-element group 196: 	39 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/req
      -- 
    req_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(196), ack => W_c4_168_delayed_14_0_177_inst_req_0); -- 
    access_T_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(76) & access_T_CP_0_elements(39) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_update_start_
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/req
      -- 
    req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(197), ack => W_c4_168_delayed_14_0_177_inst_req_1); -- 
    access_T_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	72 
    -- CP-element group 198: 	35 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/ack
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_168_delayed_14_0_177_inst_ack_0, ack => access_T_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/ack
      -- 
    ack_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_168_delayed_14_0_177_inst_ack_1, ack => access_T_CP_0_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	199 
    -- CP-element group 200: 	174 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => WPIPE_input_pipe1_181_inst_req_0); -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(195) & access_T_CP_0_elements(199) & access_T_CP_0_elements(174) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	197 
    -- CP-element group 201: 	172 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_update_start_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/req
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_181_inst_ack_0, ack => access_T_CP_0_elements(201)); -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => WPIPE_input_pipe1_181_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: 	179 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/ack
      -- 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_181_inst_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	10 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	151 
    -- CP-element group 204: 	12 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	6 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/$exit
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(202) & access_T_CP_0_elements(151) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	5 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/$exit
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/ack
      -- 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	5 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/$exit
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/ack
      -- 
    ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	3 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	1 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_26/do_while_stmt_44/$exit
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_44_terminator_636: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_44_terminator_636", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(206),loop_terminate => access_T_CP_0_elements(205),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_46_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(23);
      access_T_CP_0_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(26);
      access_T_CP_0_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(32);
      access_T_CP_0_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(33);
      access_T_CP_0_elements(22) <= phi_mux_reqs(1);
      phi_stmt_46_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_46_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(17), 
          phi_sample_ack => access_T_CP_0_elements(18), 
          phi_update_req => access_T_CP_0_elements(19), 
          phi_update_ack => access_T_CP_0_elements(20), 
          phi_mux_ack => access_T_CP_0_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_51_phi_seq_122_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(51);
      access_T_CP_0_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(52);
      access_T_CP_0_elements(41) <= phi_mux_reqs(1);
      phi_stmt_51_phi_seq_122 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_51_phi_seq_122") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(36), 
          phi_sample_ack => access_T_CP_0_elements(37), 
          phi_update_req => access_T_CP_0_elements(38), 
          phi_update_ack => access_T_CP_0_elements(39), 
          phi_mux_ack => access_T_CP_0_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_57_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(60);
      access_T_CP_0_elements(63)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(65);
      access_T_CP_0_elements(64)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(66);
      access_T_CP_0_elements(61) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(58);
      access_T_CP_0_elements(67)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(69);
      access_T_CP_0_elements(68)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(70);
      access_T_CP_0_elements(59) <= phi_mux_reqs(1);
      phi_stmt_57_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_57_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(55), 
          phi_sample_ack => access_T_CP_0_elements(56), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(57), 
          phi_mux_ack => access_T_CP_0_elements(62), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_61_phi_seq_230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(79);
      access_T_CP_0_elements(82)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(86);
      access_T_CP_0_elements(83)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(87);
      access_T_CP_0_elements(80) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(77);
      access_T_CP_0_elements(88)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(90);
      access_T_CP_0_elements(89)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(91);
      access_T_CP_0_elements(78) <= phi_mux_reqs(1);
      phi_stmt_61_phi_seq_230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_61_phi_seq_230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(73), 
          phi_sample_ack => access_T_CP_0_elements(74), 
          phi_update_req => access_T_CP_0_elements(75), 
          phi_update_ack => access_T_CP_0_elements(76), 
          phi_mux_ack => access_T_CP_0_elements(81), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_66_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(98);
      access_T_CP_0_elements(103)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(105);
      access_T_CP_0_elements(104)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(106);
      access_T_CP_0_elements(99) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(100);
      access_T_CP_0_elements(107)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(107);
      access_T_CP_0_elements(108)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(109);
      access_T_CP_0_elements(101) <= phi_mux_reqs(1);
      phi_stmt_66_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_66_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(94), 
          phi_sample_ack => access_T_CP_0_elements(95), 
          phi_update_req => access_T_CP_0_elements(96), 
          phi_update_ack => access_T_CP_0_elements(97), 
          phi_mux_ack => access_T_CP_0_elements(102), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_71_phi_seq_318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(121)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(123);
      access_T_CP_0_elements(122)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(124);
      access_T_CP_0_elements(117) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(118);
      access_T_CP_0_elements(125)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(125);
      access_T_CP_0_elements(126)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(119) <= phi_mux_reqs(1);
      phi_stmt_71_phi_seq_318 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_71_phi_seq_318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(113), 
          phi_update_req => access_T_CP_0_elements(114), 
          phi_update_ack => access_T_CP_0_elements(115), 
          phi_mux_ack => access_T_CP_0_elements(120), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_76_phi_seq_362_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(140)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(142);
      access_T_CP_0_elements(141)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(143);
      access_T_CP_0_elements(136) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(144)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(144);
      access_T_CP_0_elements(145)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(138) <= phi_mux_reqs(1);
      phi_stmt_76_phi_seq_362 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_76_phi_seq_362") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(131), 
          phi_sample_ack => access_T_CP_0_elements(132), 
          phi_update_req => access_T_CP_0_elements(133), 
          phi_update_ack => access_T_CP_0_elements(134), 
          phi_mux_ack => access_T_CP_0_elements(139), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_125_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_205_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_218_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_231_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_241_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_293_wire : std_logic_vector(15 downto 0);
    signal ADD_u64_u64_278_wire : std_logic_vector(63 downto 0);
    signal AND_u1_u1_107_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_114_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_213_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_227_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_228_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_94_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_260_wire : std_logic_vector(31 downto 0);
    signal EQ_u2_u1_103_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_110_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_117_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_90_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_97_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_274_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_240_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_242_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_30_wire : std_logic_vector(15 downto 0);
    signal MUL_u32_u32_249_wire : std_logic_vector(31 downto 0);
    signal MUX_206_wire : std_logic_vector(15 downto 0);
    signal MUX_219_wire : std_logic_vector(15 downto 0);
    signal MUX_300_wire : std_logic_vector(15 downto 0);
    signal MUX_306_wire : std_logic_vector(15 downto 0);
    signal NEQ_u16_u1_312_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_118_wire : std_logic_vector(0 downto 0);
    signal R_address_132_resized : std_logic_vector(13 downto 0);
    signal R_address_132_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_286_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_298_wire : std_logic_vector(15 downto 0);
    signal UGT_u16_u1_106_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_113_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_295_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_93_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_303_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_39_wire : std_logic_vector(0 downto 0);
    signal address_46 : std_logic_vector(63 downto 0);
    signal array_obj_ref_133_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_root_address : std_logic_vector(13 downto 0);
    signal c1_156_delayed_14_0_158 : std_logic_vector(0 downto 0);
    signal c1_86 : std_logic_vector(0 downto 0);
    signal c2_160_delayed_14_0_165 : std_logic_vector(0 downto 0);
    signal c2_99 : std_logic_vector(0 downto 0);
    signal c3_120 : std_logic_vector(0 downto 0);
    signal c3_164_delayed_14_0_172 : std_logic_vector(0 downto 0);
    signal c4_128 : std_logic_vector(0 downto 0);
    signal c4_168_delayed_14_0_179 : std_logic_vector(0 downto 0);
    signal col_71 : std_logic_vector(15 downto 0);
    signal col_done_198 : std_logic_vector(0 downto 0);
    signal fetch_addr_135 : std_logic_vector(31 downto 0);
    signal flag1_188 : std_logic_vector(0 downto 0);
    signal fn_blk_43 : std_logic_vector(15 downto 0);
    signal konst_102_wire_constant : std_logic_vector(1 downto 0);
    signal konst_105_wire_constant : std_logic_vector(15 downto 0);
    signal konst_109_wire_constant : std_logic_vector(1 downto 0);
    signal konst_112_wire_constant : std_logic_vector(15 downto 0);
    signal konst_116_wire_constant : std_logic_vector(1 downto 0);
    signal konst_126_wire_constant : std_logic_vector(15 downto 0);
    signal konst_202_wire_constant : std_logic_vector(15 downto 0);
    signal konst_204_wire_constant : std_logic_vector(15 downto 0);
    signal konst_215_wire_constant : std_logic_vector(15 downto 0);
    signal konst_217_wire_constant : std_logic_vector(15 downto 0);
    signal konst_230_wire_constant : std_logic_vector(15 downto 0);
    signal konst_259_wire_constant : std_logic_vector(31 downto 0);
    signal konst_267_wire_constant : std_logic_vector(1 downto 0);
    signal konst_273_wire_constant : std_logic_vector(31 downto 0);
    signal konst_277_wire_constant : std_logic_vector(63 downto 0);
    signal konst_294_wire_constant : std_logic_vector(15 downto 0);
    signal konst_296_wire_constant : std_logic_vector(15 downto 0);
    signal konst_302_wire_constant : std_logic_vector(15 downto 0);
    signal konst_305_wire_constant : std_logic_vector(15 downto 0);
    signal konst_38_wire_constant : std_logic_vector(15 downto 0);
    signal konst_41_wire_constant : std_logic_vector(15 downto 0);
    signal konst_84_wire_constant : std_logic_vector(1 downto 0);
    signal konst_89_wire_constant : std_logic_vector(1 downto 0);
    signal konst_92_wire_constant : std_logic_vector(15 downto 0);
    signal konst_96_wire_constant : std_logic_vector(1 downto 0);
    signal m_factor_32 : std_logic_vector(31 downto 0);
    signal n_address_280 : std_logic_vector(63 downto 0);
    signal n_address_280_50_buffered : std_logic_vector(63 downto 0);
    signal n_blk_308 : std_logic_vector(15 downto 0);
    signal n_blk_308_65_buffered : std_logic_vector(15 downto 0);
    signal n_col_222 : std_logic_vector(15 downto 0);
    signal n_col_222_73_buffered : std_logic_vector(15 downto 0);
    signal n_left_288 : std_logic_vector(15 downto 0);
    signal n_left_288_60_buffered : std_logic_vector(15 downto 0);
    signal n_row_234 : std_logic_vector(15 downto 0);
    signal n_row_234_78_buffered : std_logic_vector(15 downto 0);
    signal n_winr_209 : std_logic_vector(15 downto 0);
    signal n_winr_209_68_buffered : std_logic_vector(15 downto 0);
    signal n_word_start_269 : std_logic_vector(1 downto 0);
    signal n_word_start_269_56_buffered : std_logic_vector(1 downto 0);
    signal na1_244 : std_logic_vector(31 downto 0);
    signal na2_251 : std_logic_vector(31 downto 0);
    signal na3_256 : std_logic_vector(31 downto 0);
    signal na4_262 : std_logic_vector(15 downto 0);
    signal nl_start_35 : std_logic_vector(15 downto 0);
    signal nl_start_35_59_buffered : std_logic_vector(15 downto 0);
    signal num_blk_61 : std_logic_vector(15 downto 0);
    signal num_left_57 : std_logic_vector(15 downto 0);
    signal ptr_deref_138_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_138_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_76 : std_logic_vector(15 downto 0);
    signal type_cast_124_wire : std_logic_vector(15 downto 0);
    signal type_cast_248_wire : std_logic_vector(31 downto 0);
    signal type_cast_266_wire : std_logic_vector(1 downto 0);
    signal type_cast_275_wire : std_logic_vector(63 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_55_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_64_wire : std_logic_vector(15 downto 0);
    signal type_cast_70_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_75_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_80_wire_constant : std_logic_vector(15 downto 0);
    signal w1_143 : std_logic_vector(15 downto 0);
    signal w2_147 : std_logic_vector(15 downto 0);
    signal w3_151 : std_logic_vector(15 downto 0);
    signal w4_155 : std_logic_vector(15 downto 0);
    signal winr_66 : std_logic_vector(15 downto 0);
    signal winr_done_193 : std_logic_vector(0 downto 0);
    signal word_read_139 : std_logic_vector(63 downto 0);
    signal word_start_51 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_133_constant_part_of_offset <= "00000000000000";
    array_obj_ref_133_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_133_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_133_resized_base_address <= "00000000000000";
    konst_102_wire_constant <= "00";
    konst_105_wire_constant <= "0000000000000010";
    konst_109_wire_constant <= "01";
    konst_112_wire_constant <= "0000000000000001";
    konst_116_wire_constant <= "10";
    konst_126_wire_constant <= "0000000000000011";
    konst_202_wire_constant <= "0000000000000000";
    konst_204_wire_constant <= "0000000000000001";
    konst_215_wire_constant <= "0000000000000000";
    konst_217_wire_constant <= "0000000000000001";
    konst_230_wire_constant <= "0000000000000001";
    konst_259_wire_constant <= "00000000000000000000000000000011";
    konst_267_wire_constant <= "00";
    konst_273_wire_constant <= "00000000000000000000000000000010";
    konst_277_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_294_wire_constant <= "0000000000000100";
    konst_296_wire_constant <= "0000000000000100";
    konst_302_wire_constant <= "0000000000000100";
    konst_305_wire_constant <= "0000000000000100";
    konst_38_wire_constant <= "0000000000000100";
    konst_41_wire_constant <= "0000000000000100";
    konst_84_wire_constant <= "00";
    konst_89_wire_constant <= "00";
    konst_92_wire_constant <= "0000000000000001";
    konst_96_wire_constant <= "01";
    ptr_deref_138_word_offset_0 <= "00000000000000";
    type_cast_49_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_55_wire_constant <= "00";
    type_cast_70_wire_constant <= "0000000000000000";
    type_cast_75_wire_constant <= "0000000000000000";
    type_cast_80_wire_constant <= "0000000000000000";
    phi_stmt_46: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_49_wire_constant & n_address_280_50_buffered;
      req <= phi_stmt_46_req_0 & phi_stmt_46_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_46",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_46_ack_0,
          idata => idata,
          odata => address_46,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_46
    phi_stmt_51: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_55_wire_constant & n_word_start_269_56_buffered;
      req <= phi_stmt_51_req_0 & phi_stmt_51_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_51",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_51_ack_0,
          idata => idata,
          odata => word_start_51,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_51
    phi_stmt_57: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nl_start_35_59_buffered & n_left_288_60_buffered;
      req <= phi_stmt_57_req_0 & phi_stmt_57_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_57",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_57_ack_0,
          idata => idata,
          odata => num_left_57,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_57
    phi_stmt_61: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_64_wire & n_blk_308_65_buffered;
      req <= phi_stmt_61_req_0 & phi_stmt_61_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_61",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_61_ack_0,
          idata => idata,
          odata => num_blk_61,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_61
    phi_stmt_66: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_winr_209_68_buffered & type_cast_70_wire_constant;
      req <= phi_stmt_66_req_0 & phi_stmt_66_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_66",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_66_ack_0,
          idata => idata,
          odata => winr_66,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_66
    phi_stmt_71: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_col_222_73_buffered & type_cast_75_wire_constant;
      req <= phi_stmt_71_req_0 & phi_stmt_71_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_71",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_71_ack_0,
          idata => idata,
          odata => col_71,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_71
    phi_stmt_76: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_row_234_78_buffered & type_cast_80_wire_constant;
      req <= phi_stmt_76_req_0 & phi_stmt_76_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_76",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_76_ack_0,
          idata => idata,
          odata => row_76,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_76
    -- flow-through select operator MUX_206_inst
    MUX_206_wire <= konst_202_wire_constant when (winr_done_193(0) /=  '0') else ADD_u16_u16_205_wire;
    -- flow-through select operator MUX_208_inst
    n_winr_209 <= MUX_206_wire when (flag1_188(0) /=  '0') else winr_66;
    -- flow-through select operator MUX_219_inst
    MUX_219_wire <= konst_215_wire_constant when (col_done_198(0) /=  '0') else ADD_u16_u16_218_wire;
    -- flow-through select operator MUX_221_inst
    n_col_222 <= MUX_219_wire when (AND_u1_u1_213_wire(0) /=  '0') else col_71;
    -- flow-through select operator MUX_233_inst
    n_row_234 <= ADD_u16_u16_231_wire when (AND_u1_u1_228_wire(0) /=  '0') else row_76;
    -- flow-through select operator MUX_268_inst
    n_word_start_269 <= type_cast_266_wire when (flag1_188(0) /=  '0') else konst_267_wire_constant;
    -- flow-through select operator MUX_279_inst
    n_address_280 <= type_cast_275_wire when (flag1_188(0) /=  '0') else ADD_u64_u64_278_wire;
    -- flow-through select operator MUX_287_inst
    n_left_288 <= nl_start_35 when (flag1_188(0) /=  '0') else SUB_u16_u16_286_wire;
    -- flow-through select operator MUX_300_inst
    MUX_300_wire <= SUB_u16_u16_298_wire when (UGT_u16_u1_295_wire(0) /=  '0') else fn_blk_43;
    -- flow-through select operator MUX_306_inst
    MUX_306_wire <= n_left_288 when (ULT_u16_u1_303_wire(0) /=  '0') else konst_305_wire_constant;
    -- flow-through select operator MUX_307_inst
    n_blk_308 <= MUX_300_wire when (flag1_188(0) /=  '0') else MUX_306_wire;
    -- flow-through select operator MUX_42_inst
    fn_blk_43 <= num_cont_buffer when (ULT_u16_u1_39_wire(0) /=  '0') else konst_41_wire_constant;
    slice_142_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_142_inst_req_0;
      slice_142_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_142_inst_req_1;
      slice_142_inst_ack_1<= update_ack(0);
      slice_142_inst: SliceSplitProtocol generic map(name => "slice_142_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w1_143, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_146_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_146_inst_req_0;
      slice_146_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_146_inst_req_1;
      slice_146_inst_ack_1<= update_ack(0);
      slice_146_inst: SliceSplitProtocol generic map(name => "slice_146_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w2_147, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_150_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_150_inst_req_0;
      slice_150_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_150_inst_req_1;
      slice_150_inst_ack_1<= update_ack(0);
      slice_150_inst: SliceSplitProtocol generic map(name => "slice_150_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w3_151, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_154_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_154_inst_req_0;
      slice_154_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_154_inst_req_1;
      slice_154_inst_ack_1<= update_ack(0);
      slice_154_inst: SliceSplitProtocol generic map(name => "slice_154_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w4_155, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_c1_156_delayed_14_0_156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c1_156_delayed_14_0_156_inst_req_0;
      W_c1_156_delayed_14_0_156_inst_ack_0<= wack(0);
      rreq(0) <= W_c1_156_delayed_14_0_156_inst_req_1;
      W_c1_156_delayed_14_0_156_inst_ack_1<= rack(0);
      W_c1_156_delayed_14_0_156_inst : InterlockBuffer generic map ( -- 
        name => "W_c1_156_delayed_14_0_156_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c1_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c1_156_delayed_14_0_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c2_160_delayed_14_0_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c2_160_delayed_14_0_163_inst_req_0;
      W_c2_160_delayed_14_0_163_inst_ack_0<= wack(0);
      rreq(0) <= W_c2_160_delayed_14_0_163_inst_req_1;
      W_c2_160_delayed_14_0_163_inst_ack_1<= rack(0);
      W_c2_160_delayed_14_0_163_inst : InterlockBuffer generic map ( -- 
        name => "W_c2_160_delayed_14_0_163_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c2_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c2_160_delayed_14_0_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c3_164_delayed_14_0_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c3_164_delayed_14_0_170_inst_req_0;
      W_c3_164_delayed_14_0_170_inst_ack_0<= wack(0);
      rreq(0) <= W_c3_164_delayed_14_0_170_inst_req_1;
      W_c3_164_delayed_14_0_170_inst_ack_1<= rack(0);
      W_c3_164_delayed_14_0_170_inst : InterlockBuffer generic map ( -- 
        name => "W_c3_164_delayed_14_0_170_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c3_120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c3_164_delayed_14_0_172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c4_168_delayed_14_0_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c4_168_delayed_14_0_177_inst_req_0;
      W_c4_168_delayed_14_0_177_inst_ack_0<= wack(0);
      rreq(0) <= W_c4_168_delayed_14_0_177_inst_req_1;
      W_c4_168_delayed_14_0_177_inst_ack_1<= rack(0);
      W_c4_168_delayed_14_0_177_inst : InterlockBuffer generic map ( -- 
        name => "W_c4_168_delayed_14_0_177_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c4_128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c4_168_delayed_14_0_179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nl_start_33_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := num_cont_buffer(15 downto 0);
      nl_start_35 <= tmp_var; -- 
    end process;
    addr_of_134_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_134_final_reg_req_0;
      addr_of_134_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_134_final_reg_req_1;
      addr_of_134_final_reg_ack_1<= rack(0);
      addr_of_134_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_134_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_133_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address_280_50_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_280_50_buf_req_0;
      n_address_280_50_buf_ack_0<= wack(0);
      rreq(0) <= n_address_280_50_buf_req_1;
      n_address_280_50_buf_ack_1<= rack(0);
      n_address_280_50_buf : InterlockBuffer generic map ( -- 
        name => "n_address_280_50_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_280_50_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_blk_308_65_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_blk_308_65_buf_req_0;
      n_blk_308_65_buf_ack_0<= wack(0);
      rreq(0) <= n_blk_308_65_buf_req_1;
      n_blk_308_65_buf_ack_1<= rack(0);
      n_blk_308_65_buf : InterlockBuffer generic map ( -- 
        name => "n_blk_308_65_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_blk_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_blk_308_65_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_222_73_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_222_73_buf_req_0;
      n_col_222_73_buf_ack_0<= wack(0);
      rreq(0) <= n_col_222_73_buf_req_1;
      n_col_222_73_buf_ack_1<= rack(0);
      n_col_222_73_buf : InterlockBuffer generic map ( -- 
        name => "n_col_222_73_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_222_73_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_left_288_60_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_left_288_60_buf_req_0;
      n_left_288_60_buf_ack_0<= wack(0);
      rreq(0) <= n_left_288_60_buf_req_1;
      n_left_288_60_buf_ack_1<= rack(0);
      n_left_288_60_buf : InterlockBuffer generic map ( -- 
        name => "n_left_288_60_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_left_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_left_288_60_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_234_78_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_234_78_buf_req_0;
      n_row_234_78_buf_ack_0<= wack(0);
      rreq(0) <= n_row_234_78_buf_req_1;
      n_row_234_78_buf_ack_1<= rack(0);
      n_row_234_78_buf : InterlockBuffer generic map ( -- 
        name => "n_row_234_78_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_234_78_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_winr_209_68_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_winr_209_68_buf_req_0;
      n_winr_209_68_buf_ack_0<= wack(0);
      rreq(0) <= n_winr_209_68_buf_req_1;
      n_winr_209_68_buf_ack_1<= rack(0);
      n_winr_209_68_buf : InterlockBuffer generic map ( -- 
        name => "n_winr_209_68_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_winr_209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_winr_209_68_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_word_start_269_56_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_word_start_269_56_buf_req_0;
      n_word_start_269_56_buf_ack_0<= wack(0);
      rreq(0) <= n_word_start_269_56_buf_req_1;
      n_word_start_269_56_buf_ack_1<= rack(0);
      n_word_start_269_56_buf : InterlockBuffer generic map ( -- 
        name => "n_word_start_269_56_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_word_start_269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_word_start_269_56_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nl_start_35_59_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nl_start_35_59_buf_req_0;
      nl_start_35_59_buf_ack_0<= wack(0);
      rreq(0) <= nl_start_35_59_buf_req_1;
      nl_start_35_59_buf_ack_1<= rack(0);
      nl_start_35_59_buf : InterlockBuffer generic map ( -- 
        name => "nl_start_35_59_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nl_start_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nl_start_35_59_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_124_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := word_start_51(1 downto 0);
      type_cast_124_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_243_inst
    process(MUL_u16_u16_242_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_242_wire(15 downto 0);
      na1_244 <= tmp_var; -- 
    end process;
    -- interlock type_cast_248_inst
    process(n_winr_209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_winr_209(15 downto 0);
      type_cast_248_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_250_inst
    process(MUL_u32_u32_249_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := MUL_u32_u32_249_wire(31 downto 0);
      na2_251 <= tmp_var; -- 
    end process;
    -- interlock type_cast_261_inst
    process(AND_u32_u32_260_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := AND_u32_u32_260_wire(15 downto 0);
      na4_262 <= tmp_var; -- 
    end process;
    -- interlock type_cast_266_inst
    process(na4_262) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := na4_262(1 downto 0);
      type_cast_266_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_275_inst
    process(LSHR_u32_u32_274_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_274_wire(31 downto 0);
      type_cast_275_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_31_inst
    process(MUL_u16_u16_30_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_30_wire(15 downto 0);
      m_factor_32 <= tmp_var; -- 
    end process;
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_blk_43,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_64_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_133_index_1_rename
    process(R_address_132_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_132_resized;
      ov(13 downto 0) := iv;
      R_address_132_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_133_index_1_resize
    process(address_46) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_46;
      ov := iv(13 downto 0);
      R_address_132_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_133_root_address_inst
    process(array_obj_ref_133_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_133_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_133_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_addr_0
    process(ptr_deref_138_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_base_resize
    process(fetch_addr_135) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_135;
      ov := iv(13 downto 0);
      ptr_deref_138_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_gather_scatter
    process(ptr_deref_138_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_data_0;
      ov(63 downto 0) := iv;
      word_read_139 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_root_address_inst
    process(ptr_deref_138_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_44_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u16_u1_312_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_44_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_44_branch_req_0,
          ack0 => do_while_stmt_44_branch_ack_0,
          ack1 => do_while_stmt_44_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_125_inst
    process(num_blk_61, type_cast_124_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_blk_61, type_cast_124_wire, tmp_var);
      ADD_u16_u16_125_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_205_inst
    process(winr_66) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(winr_66, konst_204_wire_constant, tmp_var);
      ADD_u16_u16_205_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_218_inst
    process(col_71) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_71, konst_217_wire_constant, tmp_var);
      ADD_u16_u16_218_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_231_inst
    process(row_76) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_76, konst_230_wire_constant, tmp_var);
      ADD_u16_u16_231_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_241_inst
    process(n_col_222, MUL_u16_u16_240_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(n_col_222, MUL_u16_u16_240_wire, tmp_var);
      ADD_u16_u16_241_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_293_inst
    process(fn_blk_43, na4_262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(fn_blk_43, na4_262, tmp_var);
      ADD_u16_u16_293_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_255_inst
    process(na1_244, na2_251) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(na1_244, na2_251, tmp_var);
      na3_256 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_278_inst
    process(address_46) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_46, konst_277_wire_constant, tmp_var);
      ADD_u64_u64_278_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_107_inst
    process(EQ_u2_u1_103_wire, UGT_u16_u1_106_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_103_wire, UGT_u16_u1_106_wire, tmp_var);
      AND_u1_u1_107_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_114_inst
    process(EQ_u2_u1_110_wire, UGT_u16_u1_113_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_110_wire, UGT_u16_u1_113_wire, tmp_var);
      AND_u1_u1_114_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_213_inst
    process(winr_done_193, flag1_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_193, flag1_188, tmp_var);
      AND_u1_u1_213_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_227_inst
    process(col_done_198, flag1_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_198, flag1_188, tmp_var);
      AND_u1_u1_227_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_228_inst
    process(winr_done_193, AND_u1_u1_227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_193, AND_u1_u1_227_wire, tmp_var);
      AND_u1_u1_228_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_94_inst
    process(EQ_u2_u1_90_wire, UGT_u16_u1_93_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_90_wire, UGT_u16_u1_93_wire, tmp_var);
      AND_u1_u1_94_wire <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_260_inst
    process(na3_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(na3_256, konst_259_wire_constant, tmp_var);
      AND_u32_u32_260_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_187_inst
    process(num_left_57, num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_left_57, num_blk_61, tmp_var);
      flag1_188 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_192_inst
    process(winr_66, rk1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(winr_66, rk1_buffer, tmp_var);
      winr_done_193 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_197_inst
    process(col_71, col1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_71, col1_buffer, tmp_var);
      col_done_198 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_103_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_102_wire_constant, tmp_var);
      EQ_u2_u1_103_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_110_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_109_wire_constant, tmp_var);
      EQ_u2_u1_110_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_117_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_116_wire_constant, tmp_var);
      EQ_u2_u1_117_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_85_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_84_wire_constant, tmp_var);
      c1_86 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_90_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_89_wire_constant, tmp_var);
      EQ_u2_u1_90_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_97_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_96_wire_constant, tmp_var);
      EQ_u2_u1_97_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_274_inst
    process(na3_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(na3_256, konst_273_wire_constant, tmp_var);
      LSHR_u32_u32_274_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_240_inst
    process(ct_buffer, n_row_234) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, n_row_234, tmp_var);
      MUL_u16_u16_240_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_242_inst
    process(chl_in_buffer, ADD_u16_u16_241_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_in_buffer, ADD_u16_u16_241_wire, tmp_var);
      MUL_u16_u16_242_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_30_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_30_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_249_inst
    process(m_factor_32, type_cast_248_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(m_factor_32, type_cast_248_wire, tmp_var);
      MUL_u32_u32_249_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u16_u1_312_inst
    process(n_row_234, row1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(n_row_234, row1_buffer, tmp_var);
      NEQ_u16_u1_312_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_118_inst
    process(AND_u1_u1_114_wire, EQ_u2_u1_117_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_114_wire, EQ_u2_u1_117_wire, tmp_var);
      OR_u1_u1_118_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_119_inst
    process(AND_u1_u1_107_wire, OR_u1_u1_118_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_107_wire, OR_u1_u1_118_wire, tmp_var);
      c3_120 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_98_inst
    process(AND_u1_u1_94_wire, EQ_u2_u1_97_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_94_wire, EQ_u2_u1_97_wire, tmp_var);
      c2_99 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_286_inst
    process(num_left_57, num_blk_61) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(num_left_57, num_blk_61, tmp_var);
      SUB_u16_u16_286_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_298_inst
    process(konst_296_wire_constant, na4_262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_296_wire_constant, na4_262, tmp_var);
      SUB_u16_u16_298_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_106_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_105_wire_constant, tmp_var);
      UGT_u16_u1_106_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_113_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_112_wire_constant, tmp_var);
      UGT_u16_u1_113_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_127_inst
    process(ADD_u16_u16_125_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_125_wire, konst_126_wire_constant, tmp_var);
      c4_128 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_295_inst
    process(ADD_u16_u16_293_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_293_wire, konst_294_wire_constant, tmp_var);
      UGT_u16_u1_295_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_93_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_92_wire_constant, tmp_var);
      UGT_u16_u1_93_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_303_inst
    process(n_left_288) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_left_288, konst_302_wire_constant, tmp_var);
      ULT_u16_u1_303_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_39_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(num_cont_buffer, konst_38_wire_constant, tmp_var);
      ULT_u16_u1_39_wire <= tmp_var; --
    end process;
    -- shared split operator group (42) : array_obj_ref_133_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_132_scaled;
      array_obj_ref_133_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_133_index_offset_req_0;
      array_obj_ref_133_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_133_index_offset_req_1;
      array_obj_ref_133_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared load operator group (0) : ptr_deref_138_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_138_load_0_req_0;
      ptr_deref_138_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_138_load_0_req_1;
      ptr_deref_138_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_138_word_address_0;
      ptr_deref_138_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_174_inst WPIPE_input_pipe1_167_inst WPIPE_input_pipe1_160_inst WPIPE_input_pipe1_181_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_174_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_167_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_160_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_181_inst_req_0;
      WPIPE_input_pipe1_174_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_167_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_160_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_181_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_174_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_167_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_160_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_181_inst_req_1;
      WPIPE_input_pipe1_174_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_167_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_160_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_181_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= c4_168_delayed_14_0_179(0);
      guard_vector(1)  <= c1_156_delayed_14_0_158(0);
      guard_vector(2)  <= c2_160_delayed_14_0_165(0);
      guard_vector(3)  <= c3_164_delayed_14_0_172(0);
      data_in <= w3_151 & w2_147 & w1_143 & w4_155;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(95 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1120_start: Boolean;
  signal convolution3D_CP_1120_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_500_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_524_inst_req_1 : boolean;
  signal type_cast_500_inst_ack_0 : boolean;
  signal type_cast_500_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_524_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_508_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_526_inst_req_0 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_555_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_601_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_541_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_588_inst_req_0 : boolean;
  signal type_cast_500_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_588_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_601_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_493_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_601_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_557_inst_ack_1 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_572_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_557_inst_req_1 : boolean;
  signal type_cast_577_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_541_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_588_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_493_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_526_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_493_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_603_inst_req_1 : boolean;
  signal type_cast_515_inst_req_1 : boolean;
  signal type_cast_577_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_601_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_572_inst_ack_0 : boolean;
  signal type_cast_546_inst_ack_0 : boolean;
  signal type_cast_531_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_508_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_557_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_557_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_603_inst_ack_0 : boolean;
  signal type_cast_562_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_588_inst_ack_0 : boolean;
  signal type_cast_515_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_526_inst_req_1 : boolean;
  signal type_cast_577_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_524_inst_ack_0 : boolean;
  signal type_cast_546_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_555_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_510_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_555_inst_req_1 : boolean;
  signal type_cast_484_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_510_inst_req_0 : boolean;
  signal type_cast_546_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_603_inst_req_0 : boolean;
  signal type_cast_531_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_526_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_940_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_961_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_961_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_617_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_603_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_req_0 : boolean;
  signal ptr_deref_974_store_0_req_1 : boolean;
  signal type_cast_515_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_495_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_493_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_586_inst_req_0 : boolean;
  signal type_cast_531_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_524_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_617_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_555_inst_ack_0 : boolean;
  signal type_cast_531_inst_ack_1 : boolean;
  signal type_cast_608_inst_req_0 : boolean;
  signal type_cast_562_inst_ack_1 : boolean;
  signal type_cast_515_inst_ack_1 : boolean;
  signal type_cast_562_inst_req_0 : boolean;
  signal type_cast_484_inst_ack_1 : boolean;
  signal type_cast_546_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_req_1 : boolean;
  signal type_cast_562_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_572_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_572_inst_ack_1 : boolean;
  signal type_cast_593_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_539_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_495_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_586_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_617_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_619_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_617_inst_req_0 : boolean;
  signal type_cast_624_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1088_inst_ack_1 : boolean;
  signal type_cast_624_inst_ack_1 : boolean;
  signal type_cast_608_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1679_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_619_inst_req_0 : boolean;
  signal type_cast_1167_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_619_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_940_inst_ack_0 : boolean;
  signal type_cast_624_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_938_inst_ack_1 : boolean;
  signal type_cast_608_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_634_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_634_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1088_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_539_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_619_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_586_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_541_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_ack_1 : boolean;
  signal ptr_deref_1160_store_0_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_938_inst_req_1 : boolean;
  signal type_cast_577_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_634_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1088_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_634_inst_ack_1 : boolean;
  signal ptr_deref_1160_store_0_req_1 : boolean;
  signal type_cast_624_inst_req_0 : boolean;
  signal type_cast_608_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_539_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_508_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_495_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_586_inst_req_1 : boolean;
  signal type_cast_593_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_940_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_495_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_510_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_510_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_541_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_508_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_539_inst_ack_0 : boolean;
  signal type_cast_1167_inst_req_1 : boolean;
  signal type_cast_966_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_961_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_437_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_437_inst_ack_0 : boolean;
  signal ptr_deref_974_store_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_437_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_437_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_441_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_441_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_441_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_441_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_446_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_446_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_446_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_961_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_446_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_448_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_448_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_448_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_448_inst_ack_1 : boolean;
  signal type_cast_453_inst_req_0 : boolean;
  signal type_cast_453_inst_ack_0 : boolean;
  signal type_cast_453_inst_req_1 : boolean;
  signal type_cast_453_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_462_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_462_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_462_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_462_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_464_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_464_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_464_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_464_inst_ack_1 : boolean;
  signal type_cast_469_inst_req_0 : boolean;
  signal type_cast_469_inst_ack_0 : boolean;
  signal type_cast_469_inst_req_1 : boolean;
  signal type_cast_469_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_477_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_477_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_477_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_477_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_479_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_479_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_479_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_479_inst_ack_1 : boolean;
  signal type_cast_484_inst_req_0 : boolean;
  signal type_cast_484_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1088_inst_req_0 : boolean;
  signal type_cast_1095_inst_ack_1 : boolean;
  signal if_stmt_1117_branch_ack_0 : boolean;
  signal type_cast_639_inst_req_0 : boolean;
  signal type_cast_639_inst_ack_0 : boolean;
  signal type_cast_639_inst_req_1 : boolean;
  signal type_cast_639_inst_ack_1 : boolean;
  signal type_cast_1167_inst_ack_0 : boolean;
  signal type_cast_1167_inst_req_0 : boolean;
  signal type_cast_1095_inst_req_1 : boolean;
  signal if_stmt_1117_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_648_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_648_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_648_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_648_inst_ack_1 : boolean;
  signal if_stmt_1117_branch_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_650_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_650_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_940_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_650_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_650_inst_ack_1 : boolean;
  signal ptr_deref_974_store_0_ack_0 : boolean;
  signal ptr_deref_974_store_0_req_0 : boolean;
  signal type_cast_655_inst_req_0 : boolean;
  signal type_cast_655_inst_ack_0 : boolean;
  signal type_cast_655_inst_req_1 : boolean;
  signal type_cast_655_inst_ack_1 : boolean;
  signal type_cast_1095_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_663_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_663_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_663_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_663_inst_ack_1 : boolean;
  signal type_cast_1110_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_665_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_665_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_959_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_665_inst_req_1 : boolean;
  signal if_stmt_1039_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_665_inst_ack_1 : boolean;
  signal type_cast_670_inst_req_0 : boolean;
  signal type_cast_670_inst_ack_0 : boolean;
  signal type_cast_670_inst_req_1 : boolean;
  signal type_cast_670_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_959_inst_req_1 : boolean;
  signal type_cast_1095_inst_req_0 : boolean;
  signal type_cast_1110_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_679_inst_req_0 : boolean;
  signal if_stmt_1039_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_679_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_938_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_679_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_679_inst_ack_1 : boolean;
  signal ptr_deref_1160_store_0_ack_0 : boolean;
  signal ptr_deref_1160_store_0_req_0 : boolean;
  signal type_cast_1110_inst_ack_0 : boolean;
  signal type_cast_1110_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_681_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_681_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_959_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_681_inst_req_1 : boolean;
  signal if_stmt_1039_branch_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_681_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_959_inst_req_0 : boolean;
  signal type_cast_686_inst_req_0 : boolean;
  signal type_cast_686_inst_ack_0 : boolean;
  signal type_cast_686_inst_req_1 : boolean;
  signal type_cast_686_inst_ack_1 : boolean;
  signal addr_of_1157_final_reg_ack_1 : boolean;
  signal type_cast_695_inst_req_0 : boolean;
  signal type_cast_695_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_938_inst_req_0 : boolean;
  signal addr_of_1157_final_reg_req_1 : boolean;
  signal type_cast_695_inst_req_1 : boolean;
  signal type_cast_695_inst_ack_1 : boolean;
  signal type_cast_699_inst_req_0 : boolean;
  signal type_cast_699_inst_ack_0 : boolean;
  signal type_cast_699_inst_req_1 : boolean;
  signal type_cast_699_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1090_inst_ack_1 : boolean;
  signal addr_of_1157_final_reg_ack_0 : boolean;
  signal type_cast_715_inst_req_0 : boolean;
  signal if_stmt_988_branch_ack_0 : boolean;
  signal type_cast_715_inst_ack_0 : boolean;
  signal addr_of_1157_final_reg_req_0 : boolean;
  signal type_cast_715_inst_req_1 : boolean;
  signal type_cast_715_inst_ack_1 : boolean;
  signal type_cast_945_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1090_inst_req_1 : boolean;
  signal type_cast_945_inst_req_1 : boolean;
  signal array_obj_ref_1156_index_offset_ack_1 : boolean;
  signal array_obj_ref_1156_index_offset_req_1 : boolean;
  signal array_obj_ref_1156_index_offset_ack_0 : boolean;
  signal array_obj_ref_1156_index_offset_req_0 : boolean;
  signal if_stmt_723_branch_req_0 : boolean;
  signal if_stmt_723_branch_ack_1 : boolean;
  signal if_stmt_723_branch_ack_0 : boolean;
  signal type_cast_743_inst_req_0 : boolean;
  signal if_stmt_988_branch_ack_1 : boolean;
  signal type_cast_743_inst_ack_0 : boolean;
  signal type_cast_743_inst_req_1 : boolean;
  signal type_cast_743_inst_ack_1 : boolean;
  signal type_cast_945_inst_ack_0 : boolean;
  signal type_cast_966_inst_ack_1 : boolean;
  signal type_cast_966_inst_req_1 : boolean;
  signal type_cast_759_inst_req_0 : boolean;
  signal type_cast_759_inst_ack_0 : boolean;
  signal type_cast_759_inst_req_1 : boolean;
  signal if_stmt_988_branch_req_0 : boolean;
  signal type_cast_759_inst_ack_1 : boolean;
  signal type_cast_945_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1090_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1090_inst_req_0 : boolean;
  signal type_cast_966_inst_ack_0 : boolean;
  signal type_cast_768_inst_req_0 : boolean;
  signal type_cast_768_inst_ack_0 : boolean;
  signal type_cast_768_inst_req_1 : boolean;
  signal type_cast_768_inst_ack_1 : boolean;
  signal type_cast_778_inst_req_0 : boolean;
  signal type_cast_778_inst_ack_0 : boolean;
  signal ptr_deref_1470_store_0_req_0 : boolean;
  signal type_cast_778_inst_req_1 : boolean;
  signal type_cast_778_inst_ack_1 : boolean;
  signal ptr_deref_1470_store_0_ack_0 : boolean;
  signal array_obj_ref_813_index_offset_req_0 : boolean;
  signal array_obj_ref_813_index_offset_ack_0 : boolean;
  signal array_obj_ref_813_index_offset_req_1 : boolean;
  signal array_obj_ref_813_index_offset_ack_1 : boolean;
  signal type_cast_1610_inst_req_0 : boolean;
  signal if_stmt_1484_branch_ack_1 : boolean;
  signal addr_of_814_final_reg_req_0 : boolean;
  signal addr_of_814_final_reg_ack_0 : boolean;
  signal addr_of_814_final_reg_req_1 : boolean;
  signal addr_of_814_final_reg_ack_1 : boolean;
  signal type_cast_1550_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_817_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_817_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_817_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_817_inst_ack_1 : boolean;
  signal type_cast_1610_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_819_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_819_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_819_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_819_inst_ack_1 : boolean;
  signal type_cast_1610_inst_req_1 : boolean;
  signal type_cast_1758_inst_ack_1 : boolean;
  signal type_cast_824_inst_req_0 : boolean;
  signal type_cast_824_inst_ack_0 : boolean;
  signal type_cast_824_inst_req_1 : boolean;
  signal type_cast_1610_inst_ack_1 : boolean;
  signal type_cast_824_inst_ack_1 : boolean;
  signal type_cast_1758_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_833_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_833_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_833_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_833_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_835_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_835_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_835_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_835_inst_ack_1 : boolean;
  signal if_stmt_1617_branch_req_0 : boolean;
  signal type_cast_1710_inst_req_0 : boolean;
  signal type_cast_840_inst_req_0 : boolean;
  signal type_cast_840_inst_ack_0 : boolean;
  signal type_cast_1710_inst_ack_0 : boolean;
  signal type_cast_840_inst_req_1 : boolean;
  signal type_cast_840_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_854_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_854_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_854_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_854_inst_ack_1 : boolean;
  signal if_stmt_1617_branch_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_856_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_856_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_856_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_856_inst_ack_1 : boolean;
  signal type_cast_861_inst_req_0 : boolean;
  signal type_cast_861_inst_ack_0 : boolean;
  signal type_cast_861_inst_req_1 : boolean;
  signal type_cast_861_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_875_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_875_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_875_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_875_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_877_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_877_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_877_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_877_inst_ack_1 : boolean;
  signal type_cast_882_inst_req_0 : boolean;
  signal type_cast_882_inst_ack_0 : boolean;
  signal type_cast_882_inst_req_1 : boolean;
  signal type_cast_882_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_896_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_896_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_896_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_896_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_898_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_898_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_898_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_898_inst_ack_1 : boolean;
  signal type_cast_903_inst_req_0 : boolean;
  signal type_cast_903_inst_ack_0 : boolean;
  signal type_cast_903_inst_req_1 : boolean;
  signal type_cast_903_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_917_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_917_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_917_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_917_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_919_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_919_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_919_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_919_inst_ack_1 : boolean;
  signal type_cast_924_inst_req_0 : boolean;
  signal type_cast_924_inst_ack_0 : boolean;
  signal type_cast_924_inst_req_1 : boolean;
  signal type_cast_924_inst_ack_1 : boolean;
  signal type_cast_1171_inst_req_0 : boolean;
  signal type_cast_1171_inst_ack_0 : boolean;
  signal type_cast_1171_inst_req_1 : boolean;
  signal type_cast_1171_inst_ack_1 : boolean;
  signal type_cast_1175_inst_req_0 : boolean;
  signal type_cast_1175_inst_ack_0 : boolean;
  signal type_cast_1175_inst_req_1 : boolean;
  signal type_cast_1175_inst_ack_1 : boolean;
  signal type_cast_1762_inst_req_0 : boolean;
  signal ptr_deref_1660_store_0_ack_1 : boolean;
  signal type_cast_1595_inst_ack_1 : boolean;
  signal ptr_deref_1660_store_0_req_1 : boolean;
  signal type_cast_1179_inst_req_0 : boolean;
  signal type_cast_1179_inst_ack_0 : boolean;
  signal type_cast_1179_inst_req_1 : boolean;
  signal type_cast_1179_inst_ack_1 : boolean;
  signal type_cast_1595_inst_req_1 : boolean;
  signal if_stmt_1484_branch_req_0 : boolean;
  signal if_stmt_1217_branch_req_0 : boolean;
  signal if_stmt_1217_branch_ack_1 : boolean;
  signal if_stmt_1617_branch_ack_0 : boolean;
  signal if_stmt_1217_branch_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1679_inst_req_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal ptr_deref_1470_store_0_ack_1 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal type_cast_1729_inst_ack_1 : boolean;
  signal type_cast_1729_inst_req_1 : boolean;
  signal type_cast_1720_inst_ack_1 : boolean;
  signal type_cast_1242_inst_req_0 : boolean;
  signal type_cast_1242_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1686_inst_ack_1 : boolean;
  signal type_cast_1242_inst_req_1 : boolean;
  signal type_cast_1242_inst_ack_1 : boolean;
  signal type_cast_1595_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1686_inst_req_1 : boolean;
  signal type_cast_1251_inst_req_0 : boolean;
  signal type_cast_1251_inst_ack_0 : boolean;
  signal type_cast_1251_inst_req_1 : boolean;
  signal addr_of_1657_final_reg_ack_1 : boolean;
  signal type_cast_1251_inst_ack_1 : boolean;
  signal type_cast_1729_inst_ack_0 : boolean;
  signal type_cast_1729_inst_req_0 : boolean;
  signal ptr_deref_1660_store_0_ack_0 : boolean;
  signal ptr_deref_1660_store_0_req_0 : boolean;
  signal type_cast_1595_inst_req_0 : boolean;
  signal type_cast_1260_inst_req_0 : boolean;
  signal addr_of_1657_final_reg_req_1 : boolean;
  signal type_cast_1260_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1686_inst_ack_0 : boolean;
  signal type_cast_1260_inst_req_1 : boolean;
  signal type_cast_1260_inst_ack_1 : boolean;
  signal type_cast_1758_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1686_inst_req_0 : boolean;
  signal type_cast_1269_inst_req_0 : boolean;
  signal addr_of_1657_final_reg_ack_0 : boolean;
  signal type_cast_1269_inst_ack_0 : boolean;
  signal type_cast_1269_inst_req_1 : boolean;
  signal addr_of_1657_final_reg_req_0 : boolean;
  signal type_cast_1269_inst_ack_1 : boolean;
  signal type_cast_1758_inst_req_0 : boolean;
  signal type_cast_1274_inst_req_0 : boolean;
  signal type_cast_1274_inst_ack_0 : boolean;
  signal type_cast_1274_inst_req_1 : boolean;
  signal type_cast_1274_inst_ack_1 : boolean;
  signal type_cast_1720_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1590_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1590_inst_req_1 : boolean;
  signal ptr_deref_1470_store_0_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1590_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1590_inst_req_0 : boolean;
  signal array_obj_ref_1309_index_offset_req_0 : boolean;
  signal array_obj_ref_1309_index_offset_ack_0 : boolean;
  signal array_obj_ref_1309_index_offset_req_1 : boolean;
  signal array_obj_ref_1309_index_offset_ack_1 : boolean;
  signal array_obj_ref_1656_index_offset_ack_1 : boolean;
  signal array_obj_ref_1656_index_offset_req_1 : boolean;
  signal addr_of_1310_final_reg_req_0 : boolean;
  signal addr_of_1310_final_reg_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1682_inst_ack_1 : boolean;
  signal addr_of_1310_final_reg_req_1 : boolean;
  signal addr_of_1310_final_reg_ack_1 : boolean;
  signal if_stmt_1535_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1313_inst_req_0 : boolean;
  signal array_obj_ref_1656_index_offset_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1313_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1313_inst_req_1 : boolean;
  signal array_obj_ref_1656_index_offset_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1313_inst_ack_1 : boolean;
  signal type_cast_1720_inst_ack_0 : boolean;
  signal type_cast_1720_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1679_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1679_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1315_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1315_inst_ack_0 : boolean;
  signal if_stmt_1535_branch_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1315_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1315_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1588_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1588_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1682_inst_req_1 : boolean;
  signal type_cast_1320_inst_req_0 : boolean;
  signal type_cast_1320_inst_ack_0 : boolean;
  signal type_cast_1320_inst_req_1 : boolean;
  signal type_cast_1320_inst_ack_1 : boolean;
  signal if_stmt_1535_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1329_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1329_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1329_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1329_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1331_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1331_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1331_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1331_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1588_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1588_inst_req_0 : boolean;
  signal type_cast_1336_inst_req_0 : boolean;
  signal type_cast_1336_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1682_inst_ack_0 : boolean;
  signal type_cast_1336_inst_req_1 : boolean;
  signal type_cast_1336_inst_ack_1 : boolean;
  signal type_cast_1762_inst_ack_0 : boolean;
  signal call_stmt_1667_call_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1350_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1350_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1350_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1350_inst_ack_1 : boolean;
  signal call_stmt_1667_call_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1352_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1352_inst_ack_0 : boolean;
  signal type_cast_1710_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1352_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1352_inst_ack_1 : boolean;
  signal type_cast_1710_inst_req_1 : boolean;
  signal type_cast_1550_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1682_inst_req_0 : boolean;
  signal type_cast_1357_inst_req_0 : boolean;
  signal type_cast_1357_inst_ack_0 : boolean;
  signal type_cast_1357_inst_req_1 : boolean;
  signal type_cast_1357_inst_ack_1 : boolean;
  signal call_stmt_1667_call_ack_0 : boolean;
  signal call_stmt_1667_call_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1371_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1371_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1371_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1371_inst_ack_1 : boolean;
  signal type_cast_1550_inst_req_1 : boolean;
  signal type_cast_1550_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1373_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1373_inst_ack_0 : boolean;
  signal if_stmt_1484_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1373_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1373_inst_ack_1 : boolean;
  signal type_cast_1378_inst_req_0 : boolean;
  signal type_cast_1378_inst_ack_0 : boolean;
  signal type_cast_1378_inst_req_1 : boolean;
  signal type_cast_1378_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1394_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1394_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1394_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1394_inst_ack_1 : boolean;
  signal type_cast_1399_inst_req_0 : boolean;
  signal type_cast_1399_inst_ack_0 : boolean;
  signal type_cast_1399_inst_req_1 : boolean;
  signal type_cast_1399_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1413_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1413_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1413_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1413_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1415_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1415_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1415_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1415_inst_ack_1 : boolean;
  signal type_cast_1420_inst_req_0 : boolean;
  signal type_cast_1420_inst_ack_0 : boolean;
  signal type_cast_1420_inst_req_1 : boolean;
  signal type_cast_1420_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1434_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1434_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1434_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1434_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1436_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1436_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1436_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1436_inst_ack_1 : boolean;
  signal type_cast_1441_inst_req_0 : boolean;
  signal type_cast_1441_inst_ack_0 : boolean;
  signal type_cast_1441_inst_req_1 : boolean;
  signal type_cast_1441_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1455_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1455_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1455_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1455_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1457_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1457_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1457_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1457_inst_ack_1 : boolean;
  signal type_cast_1462_inst_req_0 : boolean;
  signal type_cast_1462_inst_ack_0 : boolean;
  signal type_cast_1462_inst_req_1 : boolean;
  signal type_cast_1462_inst_ack_1 : boolean;
  signal type_cast_1762_inst_req_1 : boolean;
  signal type_cast_1762_inst_ack_1 : boolean;
  signal call_stmt_1766_call_req_0 : boolean;
  signal call_stmt_1766_call_ack_0 : boolean;
  signal call_stmt_1766_call_req_1 : boolean;
  signal call_stmt_1766_call_ack_1 : boolean;
  signal call_stmt_1773_call_req_0 : boolean;
  signal call_stmt_1773_call_ack_0 : boolean;
  signal call_stmt_1773_call_req_1 : boolean;
  signal call_stmt_1773_call_ack_1 : boolean;
  signal if_stmt_1785_branch_req_0 : boolean;
  signal if_stmt_1785_branch_ack_1 : boolean;
  signal if_stmt_1785_branch_ack_0 : boolean;
  signal type_cast_1795_inst_req_0 : boolean;
  signal type_cast_1795_inst_ack_0 : boolean;
  signal type_cast_1795_inst_req_1 : boolean;
  signal type_cast_1795_inst_ack_1 : boolean;
  signal call_stmt_1799_call_req_0 : boolean;
  signal call_stmt_1799_call_ack_0 : boolean;
  signal call_stmt_1799_call_req_1 : boolean;
  signal call_stmt_1799_call_ack_1 : boolean;
  signal type_cast_1803_inst_req_0 : boolean;
  signal type_cast_1803_inst_ack_0 : boolean;
  signal type_cast_1803_inst_req_1 : boolean;
  signal type_cast_1803_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1810_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1810_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1810_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1810_inst_ack_1 : boolean;
  signal phi_stmt_801_req_0 : boolean;
  signal type_cast_807_inst_req_0 : boolean;
  signal type_cast_807_inst_ack_0 : boolean;
  signal type_cast_807_inst_req_1 : boolean;
  signal type_cast_807_inst_ack_1 : boolean;
  signal phi_stmt_801_req_1 : boolean;
  signal phi_stmt_801_ack_0 : boolean;
  signal phi_stmt_1019_req_1 : boolean;
  signal type_cast_1022_inst_req_0 : boolean;
  signal type_cast_1022_inst_ack_0 : boolean;
  signal type_cast_1022_inst_req_1 : boolean;
  signal type_cast_1022_inst_ack_1 : boolean;
  signal phi_stmt_1019_req_0 : boolean;
  signal phi_stmt_1019_ack_0 : boolean;
  signal phi_stmt_1060_req_0 : boolean;
  signal phi_stmt_1067_req_0 : boolean;
  signal type_cast_1066_inst_req_0 : boolean;
  signal type_cast_1066_inst_ack_0 : boolean;
  signal type_cast_1066_inst_req_1 : boolean;
  signal type_cast_1066_inst_ack_1 : boolean;
  signal phi_stmt_1060_req_1 : boolean;
  signal type_cast_1073_inst_req_0 : boolean;
  signal type_cast_1073_inst_ack_0 : boolean;
  signal type_cast_1073_inst_req_1 : boolean;
  signal type_cast_1073_inst_ack_1 : boolean;
  signal phi_stmt_1067_req_1 : boolean;
  signal phi_stmt_1060_ack_0 : boolean;
  signal phi_stmt_1067_ack_0 : boolean;
  signal type_cast_1127_inst_req_0 : boolean;
  signal type_cast_1127_inst_ack_0 : boolean;
  signal type_cast_1127_inst_req_1 : boolean;
  signal type_cast_1127_inst_ack_1 : boolean;
  signal phi_stmt_1124_req_0 : boolean;
  signal phi_stmt_1124_ack_0 : boolean;
  signal phi_stmt_1297_req_0 : boolean;
  signal type_cast_1303_inst_req_0 : boolean;
  signal type_cast_1303_inst_ack_0 : boolean;
  signal type_cast_1303_inst_req_1 : boolean;
  signal type_cast_1303_inst_ack_1 : boolean;
  signal phi_stmt_1297_req_1 : boolean;
  signal phi_stmt_1297_ack_0 : boolean;
  signal type_cast_1521_inst_req_0 : boolean;
  signal type_cast_1521_inst_ack_0 : boolean;
  signal type_cast_1521_inst_req_1 : boolean;
  signal type_cast_1521_inst_ack_1 : boolean;
  signal phi_stmt_1515_req_1 : boolean;
  signal phi_stmt_1515_req_0 : boolean;
  signal phi_stmt_1515_ack_0 : boolean;
  signal phi_stmt_1560_req_0 : boolean;
  signal phi_stmt_1567_req_0 : boolean;
  signal type_cast_1566_inst_req_0 : boolean;
  signal type_cast_1566_inst_ack_0 : boolean;
  signal type_cast_1566_inst_req_1 : boolean;
  signal type_cast_1566_inst_ack_1 : boolean;
  signal phi_stmt_1560_req_1 : boolean;
  signal type_cast_1573_inst_req_0 : boolean;
  signal type_cast_1573_inst_ack_0 : boolean;
  signal type_cast_1573_inst_req_1 : boolean;
  signal type_cast_1573_inst_ack_1 : boolean;
  signal phi_stmt_1567_req_1 : boolean;
  signal phi_stmt_1560_ack_0 : boolean;
  signal phi_stmt_1567_ack_0 : boolean;
  signal type_cast_1627_inst_req_0 : boolean;
  signal type_cast_1627_inst_ack_0 : boolean;
  signal type_cast_1627_inst_req_1 : boolean;
  signal type_cast_1627_inst_ack_1 : boolean;
  signal phi_stmt_1624_req_0 : boolean;
  signal phi_stmt_1624_ack_0 : boolean;
  signal phi_stmt_1738_req_1 : boolean;
  signal type_cast_1741_inst_req_0 : boolean;
  signal type_cast_1741_inst_ack_0 : boolean;
  signal type_cast_1741_inst_req_1 : boolean;
  signal type_cast_1741_inst_ack_1 : boolean;
  signal phi_stmt_1738_req_0 : boolean;
  signal phi_stmt_1738_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1120_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1120: Block -- control-path 
    signal convolution3D_CP_1120_elements: BooleanArray(437 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1120_elements(0) <= convolution3D_CP_1120_start;
    convolution3D_CP_1120_symbol <= convolution3D_CP_1120_elements(369);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	46 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	88 
    -- CP-element group 0: 	95 
    -- CP-element group 0: 	102 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	116 
    -- CP-element group 0: 	119 
    -- CP-element group 0: 	122 
    -- CP-element group 0: 	125 
    -- CP-element group 0:  members (68) 
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_436/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/branch_block_stmt_436__entry__
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722__entry__
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_Update/cr
      -- 
    cr_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_500_inst_req_1); -- 
    cr_1465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_515_inst_req_1); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_577_inst_req_1); -- 
    cr_1591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_562_inst_req_1); -- 
    cr_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_484_inst_req_1); -- 
    cr_1549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_546_inst_req_1); -- 
    cr_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_531_inst_req_1); -- 
    cr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_593_inst_req_1); -- 
    cr_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_624_inst_req_1); -- 
    cr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_608_inst_req_1); -- 
    req_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => WPIPE_maxpool_output_pipe_437_inst_req_0); -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => RPIPE_maxpool_input_pipe_446_inst_req_0); -- 
    cr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_453_inst_req_1); -- 
    cr_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_469_inst_req_1); -- 
    cr_1801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_639_inst_req_1); -- 
    cr_1843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_655_inst_req_1); -- 
    cr_1885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_670_inst_req_1); -- 
    cr_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_686_inst_req_1); -- 
    cr_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_695_inst_req_1); -- 
    cr_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_699_inst_req_1); -- 
    cr_1969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_715_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_update_start_
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_Sample/ack
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_Update/req
      -- 
    ack_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_437_inst_ack_0, ack => convolution3D_CP_1120_elements(1)); -- 
    req_1241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(1), ack => WPIPE_maxpool_output_pipe_437_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_437_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_Sample/req
      -- 
    ack_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_437_inst_ack_1, ack => convolution3D_CP_1120_elements(2)); -- 
    req_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => WPIPE_maxpool_output_pipe_441_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_update_start_
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_Update/req
      -- 
    ack_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_441_inst_ack_0, ack => convolution3D_CP_1120_elements(3)); -- 
    req_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(3), ack => WPIPE_maxpool_output_pipe_441_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_441_Update/ack
      -- 
    ack_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_441_inst_ack_1, ack => convolution3D_CP_1120_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_update_start_
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_Update/cr
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_446_inst_ack_0, ack => convolution3D_CP_1120_elements(5)); -- 
    cr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(5), ack => RPIPE_maxpool_input_pipe_446_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	10 
    -- CP-element group 6: 	12 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_446_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_Sample/rr
      -- 
    ca_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_446_inst_ack_1, ack => convolution3D_CP_1120_elements(6)); -- 
    rr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(6), ack => type_cast_453_inst_req_0); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(6), ack => RPIPE_maxpool_input_pipe_462_inst_req_0); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_Sample/req
      -- 
    req_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(7), ack => WPIPE_maxpool_output_pipe_448_inst_req_0); -- 
    convolution3D_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "convolution3D_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(4) & convolution3D_CP_1120_elements(6);
      gj_convolution3D_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_update_start_
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_Sample/ack
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_Update/req
      -- 
    ack_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_448_inst_ack_0, ack => convolution3D_CP_1120_elements(8)); -- 
    req_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(8), ack => WPIPE_maxpool_output_pipe_448_inst_req_1); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_448_Update/ack
      -- 
    ack_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_448_inst_ack_1, ack => convolution3D_CP_1120_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	6 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_Sample/ra
      -- 
    ra_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_453_inst_ack_0, ack => convolution3D_CP_1120_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	123 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_453_Update/ca
      -- 
    ca_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_453_inst_ack_1, ack => convolution3D_CP_1120_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	6 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_update_start_
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_Update/cr
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_462_inst_ack_0, ack => convolution3D_CP_1120_elements(12)); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(12), ack => RPIPE_maxpool_input_pipe_462_inst_req_1); -- 
    -- CP-element group 13:  fork  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	17 
    -- CP-element group 13: 	19 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_462_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_Sample/rr
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_462_inst_ack_1, ack => convolution3D_CP_1120_elements(13)); -- 
    rr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(13), ack => type_cast_469_inst_req_0); -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(13), ack => RPIPE_maxpool_input_pipe_477_inst_req_0); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_Sample/req
      -- 
    req_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(14), ack => WPIPE_maxpool_output_pipe_464_inst_req_0); -- 
    convolution3D_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(9) & convolution3D_CP_1120_elements(13);
      gj_convolution3D_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_update_start_
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_Sample/ack
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_Update/req
      -- 
    ack_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_464_inst_ack_0, ack => convolution3D_CP_1120_elements(15)); -- 
    req_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(15), ack => WPIPE_maxpool_output_pipe_464_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_464_Update/ack
      -- 
    ack_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_464_inst_ack_1, ack => convolution3D_CP_1120_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	13 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_Sample/ra
      -- 
    ra_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_469_inst_ack_0, ack => convolution3D_CP_1120_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	123 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_469_Update/ca
      -- 
    ca_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_469_inst_ack_1, ack => convolution3D_CP_1120_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_update_start_
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_Update/cr
      -- 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_477_inst_ack_0, ack => convolution3D_CP_1120_elements(19)); -- 
    cr_1353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(19), ack => RPIPE_maxpool_input_pipe_477_inst_req_1); -- 
    -- CP-element group 20:  fork  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	26 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_477_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_Sample/rr
      -- 
    ca_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_477_inst_ack_1, ack => convolution3D_CP_1120_elements(20)); -- 
    rr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(20), ack => type_cast_484_inst_req_0); -- 
    rr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(20), ack => RPIPE_maxpool_input_pipe_493_inst_req_0); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_Sample/req
      -- 
    req_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(21), ack => WPIPE_maxpool_output_pipe_479_inst_req_0); -- 
    convolution3D_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(16) & convolution3D_CP_1120_elements(20);
      gj_convolution3D_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_update_start_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_Sample/ack
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_Update/req
      -- 
    ack_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_479_inst_ack_0, ack => convolution3D_CP_1120_elements(22)); -- 
    req_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(22), ack => WPIPE_maxpool_output_pipe_479_inst_req_1); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	28 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_479_Update/ack
      -- 
    ack_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_479_inst_ack_1, ack => convolution3D_CP_1120_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_Sample/ra
      -- 
    ra_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_484_inst_ack_0, ack => convolution3D_CP_1120_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	117 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_484_update_completed_
      -- 
    ca_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_484_inst_ack_1, ack => convolution3D_CP_1120_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	20 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_update_start_
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_Sample/$exit
      -- 
    ra_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_493_inst_ack_0, ack => convolution3D_CP_1120_elements(26)); -- 
    cr_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(26), ack => RPIPE_maxpool_input_pipe_493_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	31 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_493_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_Sample/$entry
      -- 
    ca_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_493_inst_ack_1, ack => convolution3D_CP_1120_elements(27)); -- 
    rr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(27), ack => type_cast_500_inst_req_0); -- 
    rr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(27), ack => RPIPE_maxpool_input_pipe_508_inst_req_0); -- 
    -- CP-element group 28:  join  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_Sample/req
      -- 
    req_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(28), ack => WPIPE_maxpool_output_pipe_495_inst_req_0); -- 
    convolution3D_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(23) & convolution3D_CP_1120_elements(27);
      gj_convolution3D_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_update_start_
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_Sample/ack
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_Update/req
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_Update/$entry
      -- 
    ack_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_495_inst_ack_0, ack => convolution3D_CP_1120_elements(29)); -- 
    req_1409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(29), ack => WPIPE_maxpool_output_pipe_495_inst_req_1); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_Update/ack
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_495_Update/$exit
      -- 
    ack_1410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_495_inst_ack_1, ack => convolution3D_CP_1120_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	27 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_sample_completed_
      -- 
    ra_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_500_inst_ack_0, ack => convolution3D_CP_1120_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	117 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_500_update_completed_
      -- 
    ca_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_500_inst_ack_1, ack => convolution3D_CP_1120_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	27 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_update_start_
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_Sample/$exit
      -- 
    ra_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_508_inst_ack_0, ack => convolution3D_CP_1120_elements(33)); -- 
    cr_1437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(33), ack => RPIPE_maxpool_input_pipe_508_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_508_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_sample_start_
      -- 
    ca_1438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_508_inst_ack_1, ack => convolution3D_CP_1120_elements(34)); -- 
    rr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(34), ack => type_cast_515_inst_req_0); -- 
    rr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(34), ack => RPIPE_maxpool_input_pipe_524_inst_req_0); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_Sample/req
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_sample_start_
      -- 
    req_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(35), ack => WPIPE_maxpool_output_pipe_510_inst_req_0); -- 
    convolution3D_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(30) & convolution3D_CP_1120_elements(34);
      gj_convolution3D_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_update_start_
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_Update/req
      -- 
    ack_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_510_inst_ack_0, ack => convolution3D_CP_1120_elements(36)); -- 
    req_1451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(36), ack => WPIPE_maxpool_output_pipe_510_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	42 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_510_Update/ack
      -- 
    ack_1452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_510_inst_ack_1, ack => convolution3D_CP_1120_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_Sample/ra
      -- 
    ra_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_515_inst_ack_0, ack => convolution3D_CP_1120_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	120 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_515_Update/ca
      -- 
    ca_1466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_515_inst_ack_1, ack => convolution3D_CP_1120_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_Update/cr
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_Sample/ra
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_update_start_
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_sample_completed_
      -- 
    ra_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_524_inst_ack_0, ack => convolution3D_CP_1120_elements(40)); -- 
    cr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(40), ack => RPIPE_maxpool_input_pipe_524_inst_req_1); -- 
    -- CP-element group 41:  fork  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	45 
    -- CP-element group 41: 	47 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_524_update_completed_
      -- 
    ca_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_524_inst_ack_1, ack => convolution3D_CP_1120_elements(41)); -- 
    rr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(41), ack => type_cast_531_inst_req_0); -- 
    rr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(41), ack => RPIPE_maxpool_input_pipe_539_inst_req_0); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	37 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_Sample/req
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_sample_start_
      -- 
    req_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(42), ack => WPIPE_maxpool_output_pipe_526_inst_req_0); -- 
    convolution3D_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(37) & convolution3D_CP_1120_elements(41);
      gj_convolution3D_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_update_start_
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_Update/req
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_Sample/$exit
      -- 
    ack_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_526_inst_ack_0, ack => convolution3D_CP_1120_elements(43)); -- 
    req_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(43), ack => WPIPE_maxpool_output_pipe_526_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	49 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_526_Update/ack
      -- 
    ack_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_526_inst_ack_1, ack => convolution3D_CP_1120_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	41 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_sample_completed_
      -- 
    ra_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_0, ack => convolution3D_CP_1120_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	0 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	120 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_531_Update/ca
      -- 
    ca_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_1, ack => convolution3D_CP_1120_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	41 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_update_start_
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_Update/cr
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_Sample/ra
      -- 
    ra_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_539_inst_ack_0, ack => convolution3D_CP_1120_elements(47)); -- 
    cr_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(47), ack => RPIPE_maxpool_input_pipe_539_inst_req_1); -- 
    -- CP-element group 48:  fork  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	52 
    -- CP-element group 48: 	54 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_539_Update/$exit
      -- 
    ca_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_539_inst_ack_1, ack => convolution3D_CP_1120_elements(48)); -- 
    rr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(48), ack => type_cast_546_inst_req_0); -- 
    rr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(48), ack => RPIPE_maxpool_input_pipe_555_inst_req_0); -- 
    -- CP-element group 49:  join  transition  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	44 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_sample_start_
      -- 
    req_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(49), ack => WPIPE_maxpool_output_pipe_541_inst_req_0); -- 
    convolution3D_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(44) & convolution3D_CP_1120_elements(48);
      gj_convolution3D_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_update_start_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_Update/req
      -- 
    ack_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_541_inst_ack_0, ack => convolution3D_CP_1120_elements(50)); -- 
    req_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => WPIPE_maxpool_output_pipe_541_inst_req_1); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	56 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_541_Update/$exit
      -- 
    ack_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_541_inst_ack_1, ack => convolution3D_CP_1120_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	48 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_Sample/$exit
      -- 
    ra_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_546_inst_ack_0, ack => convolution3D_CP_1120_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	126 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_546_Update/ca
      -- 
    ca_1550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_546_inst_ack_1, ack => convolution3D_CP_1120_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	48 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_update_start_
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_Update/cr
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_Sample/$exit
      -- 
    ra_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_555_inst_ack_0, ack => convolution3D_CP_1120_elements(54)); -- 
    cr_1563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(54), ack => RPIPE_maxpool_input_pipe_555_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	59 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_555_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_sample_start_
      -- 
    ca_1564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_555_inst_ack_1, ack => convolution3D_CP_1120_elements(55)); -- 
    rr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(55), ack => type_cast_562_inst_req_0); -- 
    rr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(55), ack => RPIPE_maxpool_input_pipe_570_inst_req_0); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	51 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_Sample/$entry
      -- 
    req_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(56), ack => WPIPE_maxpool_output_pipe_557_inst_req_0); -- 
    convolution3D_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(51) & convolution3D_CP_1120_elements(55);
      gj_convolution3D_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_update_start_
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_Update/req
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_sample_completed_
      -- 
    ack_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_557_inst_ack_0, ack => convolution3D_CP_1120_elements(57)); -- 
    req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(57), ack => WPIPE_maxpool_output_pipe_557_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	63 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_557_update_completed_
      -- 
    ack_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_557_inst_ack_1, ack => convolution3D_CP_1120_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	55 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_Sample/ra
      -- 
    ra_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_562_inst_ack_0, ack => convolution3D_CP_1120_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	126 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_562_Update/$exit
      -- 
    ca_1592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_562_inst_ack_1, ack => convolution3D_CP_1120_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_Update/cr
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_update_start_
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_sample_completed_
      -- 
    ra_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_570_inst_ack_0, ack => convolution3D_CP_1120_elements(61)); -- 
    cr_1605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(61), ack => RPIPE_maxpool_input_pipe_570_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	66 
    -- CP-element group 62: 	68 
    -- CP-element group 62:  members (9) 
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_570_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_Sample/$entry
      -- 
    ca_1606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_570_inst_ack_1, ack => convolution3D_CP_1120_elements(62)); -- 
    rr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(62), ack => type_cast_577_inst_req_0); -- 
    rr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(62), ack => RPIPE_maxpool_input_pipe_586_inst_req_0); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	58 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_sample_start_
      -- 
    req_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(63), ack => WPIPE_maxpool_output_pipe_572_inst_req_0); -- 
    convolution3D_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(58) & convolution3D_CP_1120_elements(62);
      gj_convolution3D_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_update_start_
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_Update/req
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_sample_completed_
      -- 
    ack_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_572_inst_ack_0, ack => convolution3D_CP_1120_elements(64)); -- 
    req_1619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(64), ack => WPIPE_maxpool_output_pipe_572_inst_req_1); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	70 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_572_Update/ack
      -- 
    ack_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_572_inst_ack_1, ack => convolution3D_CP_1120_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_Sample/$exit
      -- 
    ra_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_0, ack => convolution3D_CP_1120_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	126 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_577_update_completed_
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_1, ack => convolution3D_CP_1120_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	62 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (6) 
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_update_start_
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_Sample/ra
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_Update/cr
      -- 
    ra_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_586_inst_ack_0, ack => convolution3D_CP_1120_elements(68)); -- 
    cr_1647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(68), ack => RPIPE_maxpool_input_pipe_586_inst_req_1); -- 
    -- CP-element group 69:  fork  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: 	73 
    -- CP-element group 69: 	75 
    -- CP-element group 69:  members (9) 
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_Update/ca
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_586_Update/$exit
      -- 
    ca_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_586_inst_ack_1, ack => convolution3D_CP_1120_elements(69)); -- 
    rr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(69), ack => type_cast_593_inst_req_0); -- 
    rr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(69), ack => RPIPE_maxpool_input_pipe_601_inst_req_0); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	65 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_Sample/req
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_sample_start_
      -- 
    req_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(70), ack => WPIPE_maxpool_output_pipe_588_inst_req_0); -- 
    convolution3D_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(65) & convolution3D_CP_1120_elements(69);
      gj_convolution3D_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_Update/req
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_update_start_
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_sample_completed_
      -- 
    ack_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_588_inst_ack_0, ack => convolution3D_CP_1120_elements(71)); -- 
    req_1661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(71), ack => WPIPE_maxpool_output_pipe_588_inst_req_1); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	77 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_Update/ack
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_588_update_completed_
      -- 
    ack_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_588_inst_ack_1, ack => convolution3D_CP_1120_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_sample_completed_
      -- 
    ra_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => convolution3D_CP_1120_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	126 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_593_Update/ca
      -- 
    ca_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_1, ack => convolution3D_CP_1120_elements(74)); -- 
    -- CP-element group 75:  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	69 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (6) 
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_sample_completed_
      -- 
    ra_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_601_inst_ack_0, ack => convolution3D_CP_1120_elements(75)); -- 
    cr_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => RPIPE_maxpool_input_pipe_601_inst_req_1); -- 
    -- CP-element group 76:  fork  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	80 
    -- CP-element group 76: 	82 
    -- CP-element group 76:  members (9) 
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_601_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_Sample/rr
      -- 
    ca_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_601_inst_ack_1, ack => convolution3D_CP_1120_elements(76)); -- 
    rr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(76), ack => type_cast_608_inst_req_0); -- 
    rr_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(76), ack => RPIPE_maxpool_input_pipe_617_inst_req_0); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	72 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_Sample/req
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_Sample/$entry
      -- 
    req_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(77), ack => WPIPE_maxpool_output_pipe_603_inst_req_0); -- 
    convolution3D_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(72) & convolution3D_CP_1120_elements(76);
      gj_convolution3D_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_Update/req
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_Sample/ack
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_update_start_
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_Sample/$exit
      -- 
    ack_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_603_inst_ack_0, ack => convolution3D_CP_1120_elements(78)); -- 
    req_1703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(78), ack => WPIPE_maxpool_output_pipe_603_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	84 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_Update/ack
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_603_Update/$exit
      -- 
    ack_1704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_603_inst_ack_1, ack => convolution3D_CP_1120_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	76 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_Sample/ra
      -- 
    ra_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_0, ack => convolution3D_CP_1120_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	126 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_608_Update/ca
      -- 
    ca_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_1, ack => convolution3D_CP_1120_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	76 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_update_start_
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_sample_completed_
      -- 
    ra_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_617_inst_ack_0, ack => convolution3D_CP_1120_elements(82)); -- 
    cr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(82), ack => RPIPE_maxpool_input_pipe_617_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	87 
    -- CP-element group 83: 	89 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_617_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_Sample/rr
      -- 
    ca_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_617_inst_ack_1, ack => convolution3D_CP_1120_elements(83)); -- 
    rr_1754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(83), ack => type_cast_624_inst_req_0); -- 
    rr_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(83), ack => RPIPE_maxpool_input_pipe_632_inst_req_0); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	79 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_Sample/req
      -- 
    req_1740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(84), ack => WPIPE_maxpool_output_pipe_619_inst_req_0); -- 
    convolution3D_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(79) & convolution3D_CP_1120_elements(83);
      gj_convolution3D_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_Sample/ack
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_Update/req
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_update_start_
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_Update/$entry
      -- 
    ack_1741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_619_inst_ack_0, ack => convolution3D_CP_1120_elements(85)); -- 
    req_1745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(85), ack => WPIPE_maxpool_output_pipe_619_inst_req_1); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	91 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_Update/ack
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_619_Update/$exit
      -- 
    ack_1746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_619_inst_ack_1, ack => convolution3D_CP_1120_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_Sample/$exit
      -- 
    ra_1755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_624_inst_ack_0, ack => convolution3D_CP_1120_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	0 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	126 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_624_update_completed_
      -- 
    ca_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_624_inst_ack_1, ack => convolution3D_CP_1120_elements(88)); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	83 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_update_start_
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_Update/cr
      -- 
    ra_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_632_inst_ack_0, ack => convolution3D_CP_1120_elements(89)); -- 
    cr_1773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(89), ack => RPIPE_maxpool_input_pipe_632_inst_req_1); -- 
    -- CP-element group 90:  fork  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: 	94 
    -- CP-element group 90: 	96 
    -- CP-element group 90:  members (9) 
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_632_Update/ca
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_Sample/rr
      -- 
    ca_1774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_632_inst_ack_1, ack => convolution3D_CP_1120_elements(90)); -- 
    rr_1796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(90), ack => type_cast_639_inst_req_0); -- 
    rr_1810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(90), ack => RPIPE_maxpool_input_pipe_648_inst_req_0); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	86 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_Sample/req
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_Sample/$entry
      -- 
    req_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(91), ack => WPIPE_maxpool_output_pipe_634_inst_req_0); -- 
    convolution3D_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(86) & convolution3D_CP_1120_elements(90);
      gj_convolution3D_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_Sample/ack
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_update_start_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_Update/req
      -- 
    ack_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_634_inst_ack_0, ack => convolution3D_CP_1120_elements(92)); -- 
    req_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(92), ack => WPIPE_maxpool_output_pipe_634_inst_req_1); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	98 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_634_Update/ack
      -- 
    ack_1788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_634_inst_ack_1, ack => convolution3D_CP_1120_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	90 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_Sample/ra
      -- 
    ra_1797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_0, ack => convolution3D_CP_1120_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	0 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	126 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_639_Update/ca
      -- 
    ca_1802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_1, ack => convolution3D_CP_1120_elements(95)); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	90 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_update_start_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_Update/cr
      -- 
    ra_1811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_648_inst_ack_0, ack => convolution3D_CP_1120_elements(96)); -- 
    cr_1815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(96), ack => RPIPE_maxpool_input_pipe_648_inst_req_1); -- 
    -- CP-element group 97:  fork  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	101 
    -- CP-element group 97: 	103 
    -- CP-element group 97:  members (9) 
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_648_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_Sample/rr
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_Sample/rr
      -- 
    ca_1816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_648_inst_ack_1, ack => convolution3D_CP_1120_elements(97)); -- 
    rr_1838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(97), ack => type_cast_655_inst_req_0); -- 
    rr_1852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(97), ack => RPIPE_maxpool_input_pipe_663_inst_req_0); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	93 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_Sample/req
      -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(98), ack => WPIPE_maxpool_output_pipe_650_inst_req_0); -- 
    convolution3D_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(93) & convolution3D_CP_1120_elements(97);
      gj_convolution3D_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_update_start_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_Update/req
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_650_inst_ack_0, ack => convolution3D_CP_1120_elements(99)); -- 
    req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(99), ack => WPIPE_maxpool_output_pipe_650_inst_req_1); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	105 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_650_Update/ack
      -- 
    ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_650_inst_ack_1, ack => convolution3D_CP_1120_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_Sample/ra
      -- 
    ra_1839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_655_inst_ack_0, ack => convolution3D_CP_1120_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	0 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	126 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_655_Update/ca
      -- 
    ca_1844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_655_inst_ack_1, ack => convolution3D_CP_1120_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	97 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_update_start_
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_Update/cr
      -- 
    ra_1853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_663_inst_ack_0, ack => convolution3D_CP_1120_elements(103)); -- 
    cr_1857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(103), ack => RPIPE_maxpool_input_pipe_663_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	108 
    -- CP-element group 104: 	110 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_663_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_Sample/rr
      -- 
    ca_1858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_663_inst_ack_1, ack => convolution3D_CP_1120_elements(104)); -- 
    rr_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(104), ack => type_cast_670_inst_req_0); -- 
    rr_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(104), ack => RPIPE_maxpool_input_pipe_679_inst_req_0); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	100 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_Sample/req
      -- 
    req_1866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(105), ack => WPIPE_maxpool_output_pipe_665_inst_req_0); -- 
    convolution3D_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(100) & convolution3D_CP_1120_elements(104);
      gj_convolution3D_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_update_start_
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_Sample/ack
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_Update/req
      -- 
    ack_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_665_inst_ack_0, ack => convolution3D_CP_1120_elements(106)); -- 
    req_1871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(106), ack => WPIPE_maxpool_output_pipe_665_inst_req_1); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_665_Update/ack
      -- 
    ack_1872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_665_inst_ack_1, ack => convolution3D_CP_1120_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	104 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_Sample/ra
      -- 
    ra_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_670_inst_ack_0, ack => convolution3D_CP_1120_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	126 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_670_Update/ca
      -- 
    ca_1886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_670_inst_ack_1, ack => convolution3D_CP_1120_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	104 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_update_start_
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_Update/cr
      -- 
    ra_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_679_inst_ack_0, ack => convolution3D_CP_1120_elements(110)); -- 
    cr_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(110), ack => RPIPE_maxpool_input_pipe_679_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	115 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/RPIPE_maxpool_input_pipe_679_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_Sample/rr
      -- 
    ca_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_679_inst_ack_1, ack => convolution3D_CP_1120_elements(111)); -- 
    rr_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(111), ack => type_cast_686_inst_req_0); -- 
    -- CP-element group 112:  join  transition  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_Sample/req
      -- 
    req_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(112), ack => WPIPE_maxpool_output_pipe_681_inst_req_0); -- 
    convolution3D_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(107) & convolution3D_CP_1120_elements(111);
      gj_convolution3D_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_update_start_
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_Sample/ack
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_Update/req
      -- 
    ack_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_681_inst_ack_0, ack => convolution3D_CP_1120_elements(113)); -- 
    req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(113), ack => WPIPE_maxpool_output_pipe_681_inst_req_1); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	126 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/WPIPE_maxpool_output_pipe_681_Update/ack
      -- 
    ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_681_inst_ack_1, ack => convolution3D_CP_1120_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	111 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_Sample/ra
      -- 
    ra_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_0, ack => convolution3D_CP_1120_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	0 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	126 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_686_Update/ca
      -- 
    ca_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_1, ack => convolution3D_CP_1120_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	25 
    -- CP-element group 117: 	32 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_Sample/rr
      -- 
    rr_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(117), ack => type_cast_695_inst_req_0); -- 
    convolution3D_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(25) & convolution3D_CP_1120_elements(32);
      gj_convolution3D_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_Sample/ra
      -- 
    ra_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_0, ack => convolution3D_CP_1120_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	0 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_695_Update/ca
      -- 
    ca_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_1, ack => convolution3D_CP_1120_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	39 
    -- CP-element group 120: 	46 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_Sample/rr
      -- 
    rr_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(120), ack => type_cast_699_inst_req_0); -- 
    convolution3D_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(39) & convolution3D_CP_1120_elements(46);
      gj_convolution3D_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_Sample/ra
      -- 
    ra_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_0, ack => convolution3D_CP_1120_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	0 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_699_Update/ca
      -- 
    ca_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_1, ack => convolution3D_CP_1120_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	11 
    -- CP-element group 123: 	18 
    -- CP-element group 123: 	119 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_Sample/rr
      -- 
    rr_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(123), ack => type_cast_715_inst_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(11) & convolution3D_CP_1120_elements(18) & convolution3D_CP_1120_elements(119) & convolution3D_CP_1120_elements(122);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_Sample/ra
      -- 
    ra_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_715_inst_ack_0, ack => convolution3D_CP_1120_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	0 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/type_cast_715_Update/ca
      -- 
    ca_1970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_715_inst_ack_1, ack => convolution3D_CP_1120_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	53 
    -- CP-element group 126: 	60 
    -- CP-element group 126: 	67 
    -- CP-element group 126: 	74 
    -- CP-element group 126: 	81 
    -- CP-element group 126: 	88 
    -- CP-element group 126: 	95 
    -- CP-element group 126: 	102 
    -- CP-element group 126: 	109 
    -- CP-element group 126: 	114 
    -- CP-element group 126: 	116 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722__exit__
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_723__entry__
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_722/$exit
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_723_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_723_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_723_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_723_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_436/R_cmp447_724_place
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_723_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_723_else_link/$entry
      -- 
    branch_req_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(126), ack => if_stmt_723_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(53) & convolution3D_CP_1120_elements(60) & convolution3D_CP_1120_elements(67) & convolution3D_CP_1120_elements(74) & convolution3D_CP_1120_elements(81) & convolution3D_CP_1120_elements(88) & convolution3D_CP_1120_elements(95) & convolution3D_CP_1120_elements(102) & convolution3D_CP_1120_elements(109) & convolution3D_CP_1120_elements(114) & convolution3D_CP_1120_elements(116) & convolution3D_CP_1120_elements(125);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: 	130 
    -- CP-element group 127: 	131 
    -- CP-element group 127: 	132 
    -- CP-element group 127: 	133 
    -- CP-element group 127: 	134 
    -- CP-element group 127: 	137 
    -- CP-element group 127:  members (33) 
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_729__exit__
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798__entry__
      -- CP-element group 127: 	 branch_block_stmt_436/if_stmt_723_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/if_stmt_723_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_436/entry_bbx_xnph449
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_update_start_
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_Update/cr
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_update_start_
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_Update/cr
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_update_start_
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_Update/cr
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_update_start_
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_Update/cr
      -- CP-element group 127: 	 branch_block_stmt_436/entry_bbx_xnph449_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/entry_bbx_xnph449_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_729_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_729_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_729_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_729_PhiAck/dummy
      -- 
    if_choice_transition_1983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_723_branch_ack_1, ack => convolution3D_CP_1120_elements(127)); -- 
    rr_2000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_743_inst_req_0); -- 
    cr_2005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_743_inst_req_1); -- 
    rr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_759_inst_req_0); -- 
    cr_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_759_inst_req_1); -- 
    rr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_768_inst_req_0); -- 
    cr_2033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_768_inst_req_1); -- 
    cr_2047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_778_inst_req_1); -- 
    -- CP-element group 128:  transition  place  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	376 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_436/if_stmt_723_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_436/if_stmt_723_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_436/entry_forx_xend
      -- CP-element group 128: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1019/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/$entry
      -- 
    else_choice_transition_1987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_723_branch_ack_0, ack => convolution3D_CP_1120_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_Sample/ra
      -- 
    ra_2001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_743_inst_ack_0, ack => convolution3D_CP_1120_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	127 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	138 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_743_Update/ca
      -- 
    ca_2006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_743_inst_ack_1, ack => convolution3D_CP_1120_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	127 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_Sample/ra
      -- 
    ra_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_759_inst_ack_0, ack => convolution3D_CP_1120_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	127 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	135 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_759_Update/ca
      -- 
    ca_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_759_inst_ack_1, ack => convolution3D_CP_1120_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	127 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_Sample/ra
      -- 
    ra_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_0, ack => convolution3D_CP_1120_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	127 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_768_Update/ca
      -- 
    ca_2034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_1, ack => convolution3D_CP_1120_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	132 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_Sample/rr
      -- 
    rr_2042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(135), ack => type_cast_778_inst_req_0); -- 
    convolution3D_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(132) & convolution3D_CP_1120_elements(134);
      gj_convolution3D_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_Sample/ra
      -- 
    ra_2043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_778_inst_ack_0, ack => convolution3D_CP_1120_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	127 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/type_cast_778_Update/ca
      -- 
    ca_2048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_778_inst_ack_1, ack => convolution3D_CP_1120_elements(137)); -- 
    -- CP-element group 138:  join  transition  place  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	130 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	370 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798__exit__
      -- CP-element group 138: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody
      -- CP-element group 138: 	 branch_block_stmt_436/assign_stmt_734_to_assign_stmt_798/$exit
      -- CP-element group 138: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_801/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/$entry
      -- 
    convolution3D_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(130) & convolution3D_CP_1120_elements(137);
      gj_convolution3D_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	375 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	201 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_sample_complete
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_Sample/ack
      -- 
    ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_813_index_offset_ack_0, ack => convolution3D_CP_1120_elements(139)); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	375 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (11) 
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_root_address_calculated
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_offset_calculated
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_Update/ack
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_base_plus_offset/$entry
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_base_plus_offset/$exit
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_base_plus_offset/sum_rename_req
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_base_plus_offset/sum_rename_ack
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_request/$entry
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_request/req
      -- 
    ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_813_index_offset_ack_1, ack => convolution3D_CP_1120_elements(140)); -- 
    req_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(140), ack => addr_of_814_final_reg_req_0); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_request/$exit
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_request/ack
      -- 
    ack_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_814_final_reg_ack_0, ack => convolution3D_CP_1120_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	375 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	198 
    -- CP-element group 142:  members (19) 
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_word_addrgen/root_register_ack
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_word_addrgen/root_register_req
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_word_addrgen/$exit
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_word_addrgen/$entry
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_plus_offset/sum_rename_ack
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_plus_offset/sum_rename_req
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_plus_offset/$exit
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_plus_offset/$entry
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_addr_resize/base_resize_ack
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_addr_resize/base_resize_req
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_addr_resize/$exit
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_addr_resize/$entry
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_address_resized
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_root_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_word_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_base_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_complete/$exit
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_complete/ack
      -- 
    ack_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_814_final_reg_ack_1, ack => convolution3D_CP_1120_elements(142)); -- 
    -- CP-element group 143:  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	375 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (6) 
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_update_start_
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_Update/cr
      -- 
    ra_2106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_817_inst_ack_0, ack => convolution3D_CP_1120_elements(143)); -- 
    cr_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(143), ack => RPIPE_maxpool_input_pipe_817_inst_req_1); -- 
    -- CP-element group 144:  fork  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144: 	147 
    -- CP-element group 144: 	149 
    -- CP-element group 144:  members (12) 
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_Sample/req
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_Sample/rr
      -- 
    ca_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_817_inst_ack_1, ack => convolution3D_CP_1120_elements(144)); -- 
    req_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(144), ack => WPIPE_maxpool_output_pipe_819_inst_req_0); -- 
    rr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(144), ack => type_cast_824_inst_req_0); -- 
    rr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(144), ack => RPIPE_maxpool_input_pipe_833_inst_req_0); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_update_start_
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_Sample/ack
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_Update/req
      -- 
    ack_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_819_inst_ack_0, ack => convolution3D_CP_1120_elements(145)); -- 
    req_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(145), ack => WPIPE_maxpool_output_pipe_819_inst_req_1); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	151 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_819_Update/ack
      -- 
    ack_2125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_819_inst_ack_1, ack => convolution3D_CP_1120_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	144 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_Sample/ra
      -- 
    ra_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_824_inst_ack_0, ack => convolution3D_CP_1120_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	375 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	198 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_Update/ca
      -- 
    ca_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_824_inst_ack_1, ack => convolution3D_CP_1120_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	144 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_update_start_
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_Update/cr
      -- 
    ra_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_833_inst_ack_0, ack => convolution3D_CP_1120_elements(149)); -- 
    cr_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(149), ack => RPIPE_maxpool_input_pipe_833_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	154 
    -- CP-element group 150: 	156 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_833_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_Sample/rr
      -- 
    ca_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_833_inst_ack_1, ack => convolution3D_CP_1120_elements(150)); -- 
    rr_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => type_cast_840_inst_req_0); -- 
    rr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(150), ack => RPIPE_maxpool_input_pipe_854_inst_req_0); -- 
    -- CP-element group 151:  join  transition  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	146 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_Sample/req
      -- 
    req_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(151), ack => WPIPE_maxpool_output_pipe_835_inst_req_0); -- 
    convolution3D_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(146) & convolution3D_CP_1120_elements(150);
      gj_convolution3D_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_update_start_
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_Update/req
      -- 
    ack_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_835_inst_ack_0, ack => convolution3D_CP_1120_elements(152)); -- 
    req_2166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(152), ack => WPIPE_maxpool_output_pipe_835_inst_req_1); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	158 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_835_Update/ack
      -- 
    ack_2167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_835_inst_ack_1, ack => convolution3D_CP_1120_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	150 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_Sample/ra
      -- 
    ra_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_840_inst_ack_0, ack => convolution3D_CP_1120_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	375 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	198 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_Update/ca
      -- 
    ca_2181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_840_inst_ack_1, ack => convolution3D_CP_1120_elements(155)); -- 
    -- CP-element group 156:  transition  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	150 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (6) 
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_Update/cr
      -- 
    ra_2190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_854_inst_ack_0, ack => convolution3D_CP_1120_elements(156)); -- 
    cr_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => RPIPE_maxpool_input_pipe_854_inst_req_1); -- 
    -- CP-element group 157:  fork  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: 	161 
    -- CP-element group 157: 	163 
    -- CP-element group 157:  members (9) 
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_854_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_Sample/rr
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_Sample/rr
      -- 
    ca_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_854_inst_ack_1, ack => convolution3D_CP_1120_elements(157)); -- 
    rr_2217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(157), ack => type_cast_861_inst_req_0); -- 
    rr_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(157), ack => RPIPE_maxpool_input_pipe_875_inst_req_0); -- 
    -- CP-element group 158:  join  transition  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	153 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_Sample/req
      -- 
    req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(158), ack => WPIPE_maxpool_output_pipe_856_inst_req_0); -- 
    convolution3D_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(153) & convolution3D_CP_1120_elements(157);
      gj_convolution3D_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_update_start_
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_Sample/ack
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_Update/req
      -- 
    ack_2204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_856_inst_ack_0, ack => convolution3D_CP_1120_elements(159)); -- 
    req_2208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(159), ack => WPIPE_maxpool_output_pipe_856_inst_req_1); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	165 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_856_Update/ack
      -- 
    ack_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_856_inst_ack_1, ack => convolution3D_CP_1120_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	157 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_Sample/ra
      -- 
    ra_2218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_0, ack => convolution3D_CP_1120_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	375 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	198 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_Update/ca
      -- 
    ca_2223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_1, ack => convolution3D_CP_1120_elements(162)); -- 
    -- CP-element group 163:  transition  input  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	157 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (6) 
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_update_start_
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_Sample/ra
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_Update/cr
      -- 
    ra_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_875_inst_ack_0, ack => convolution3D_CP_1120_elements(163)); -- 
    cr_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(163), ack => RPIPE_maxpool_input_pipe_875_inst_req_1); -- 
    -- CP-element group 164:  fork  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	168 
    -- CP-element group 164: 	170 
    -- CP-element group 164:  members (9) 
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_875_Update/ca
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_Sample/rr
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_Sample/rr
      -- 
    ca_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_875_inst_ack_1, ack => convolution3D_CP_1120_elements(164)); -- 
    rr_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(164), ack => type_cast_882_inst_req_0); -- 
    rr_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(164), ack => RPIPE_maxpool_input_pipe_896_inst_req_0); -- 
    -- CP-element group 165:  join  transition  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	160 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_Sample/req
      -- 
    req_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(165), ack => WPIPE_maxpool_output_pipe_877_inst_req_0); -- 
    convolution3D_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(160) & convolution3D_CP_1120_elements(164);
      gj_convolution3D_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (6) 
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_update_start_
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_Sample/ack
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_Update/req
      -- 
    ack_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_877_inst_ack_0, ack => convolution3D_CP_1120_elements(166)); -- 
    req_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(166), ack => WPIPE_maxpool_output_pipe_877_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	172 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_877_Update/ack
      -- 
    ack_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_877_inst_ack_1, ack => convolution3D_CP_1120_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	164 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_Sample/ra
      -- 
    ra_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_882_inst_ack_0, ack => convolution3D_CP_1120_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	375 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	198 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_Update/ca
      -- 
    ca_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_882_inst_ack_1, ack => convolution3D_CP_1120_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	164 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_update_start_
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_Update/cr
      -- 
    ra_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_896_inst_ack_0, ack => convolution3D_CP_1120_elements(170)); -- 
    cr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(170), ack => RPIPE_maxpool_input_pipe_896_inst_req_1); -- 
    -- CP-element group 171:  fork  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171: 	175 
    -- CP-element group 171: 	177 
    -- CP-element group 171:  members (9) 
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_896_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_Sample/rr
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_Sample/rr
      -- 
    ca_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_896_inst_ack_1, ack => convolution3D_CP_1120_elements(171)); -- 
    rr_2301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(171), ack => type_cast_903_inst_req_0); -- 
    rr_2315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(171), ack => RPIPE_maxpool_input_pipe_917_inst_req_0); -- 
    -- CP-element group 172:  join  transition  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	167 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_Sample/req
      -- 
    req_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(172), ack => WPIPE_maxpool_output_pipe_898_inst_req_0); -- 
    convolution3D_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(167) & convolution3D_CP_1120_elements(171);
      gj_convolution3D_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_update_start_
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_Sample/ack
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_Update/req
      -- 
    ack_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_898_inst_ack_0, ack => convolution3D_CP_1120_elements(173)); -- 
    req_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(173), ack => WPIPE_maxpool_output_pipe_898_inst_req_1); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	179 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_898_Update/ack
      -- 
    ack_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_898_inst_ack_1, ack => convolution3D_CP_1120_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	171 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_Sample/ra
      -- 
    ra_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_0, ack => convolution3D_CP_1120_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	375 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	198 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_Update/ca
      -- 
    ca_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_1, ack => convolution3D_CP_1120_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	171 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_update_start_
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_Update/cr
      -- 
    ra_2316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_917_inst_ack_0, ack => convolution3D_CP_1120_elements(177)); -- 
    cr_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(177), ack => RPIPE_maxpool_input_pipe_917_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	182 
    -- CP-element group 178: 	184 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_917_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_sample_start_
      -- 
    ca_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_917_inst_ack_1, ack => convolution3D_CP_1120_elements(178)); -- 
    rr_2343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(178), ack => type_cast_924_inst_req_0); -- 
    rr_2357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(178), ack => RPIPE_maxpool_input_pipe_938_inst_req_0); -- 
    -- CP-element group 179:  join  transition  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	174 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_Sample/req
      -- 
    req_2329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(179), ack => WPIPE_maxpool_output_pipe_919_inst_req_0); -- 
    convolution3D_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(174) & convolution3D_CP_1120_elements(178);
      gj_convolution3D_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_update_start_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_Update/req
      -- 
    ack_2330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_919_inst_ack_0, ack => convolution3D_CP_1120_elements(180)); -- 
    req_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(180), ack => WPIPE_maxpool_output_pipe_919_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_919_Update/ack
      -- 
    ack_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_919_inst_ack_1, ack => convolution3D_CP_1120_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	178 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_Sample/ra
      -- 
    ra_2344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_0, ack => convolution3D_CP_1120_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	375 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	198 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_Update/ca
      -- 
    ca_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_1, ack => convolution3D_CP_1120_elements(183)); -- 
    -- CP-element group 184:  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	178 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (6) 
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_Sample/ra
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_update_start_
      -- 
    ra_2358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_938_inst_ack_0, ack => convolution3D_CP_1120_elements(184)); -- 
    cr_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(184), ack => RPIPE_maxpool_input_pipe_938_inst_req_1); -- 
    -- CP-element group 185:  fork  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185: 	189 
    -- CP-element group 185: 	191 
    -- CP-element group 185:  members (9) 
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_Sample/rr
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_938_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_Sample/rr
      -- 
    ca_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_938_inst_ack_1, ack => convolution3D_CP_1120_elements(185)); -- 
    rr_2385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(185), ack => type_cast_945_inst_req_0); -- 
    rr_2399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(185), ack => RPIPE_maxpool_input_pipe_959_inst_req_0); -- 
    -- CP-element group 186:  join  transition  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	181 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_Sample/req
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_Sample/$entry
      -- 
    req_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(186), ack => WPIPE_maxpool_output_pipe_940_inst_req_0); -- 
    convolution3D_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(181) & convolution3D_CP_1120_elements(185);
      gj_convolution3D_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_Update/req
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_update_start_
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_Sample/$exit
      -- 
    ack_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_940_inst_ack_0, ack => convolution3D_CP_1120_elements(187)); -- 
    req_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => WPIPE_maxpool_output_pipe_940_inst_req_1); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_940_update_completed_
      -- 
    ack_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_940_inst_ack_1, ack => convolution3D_CP_1120_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	185 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_Sample/$exit
      -- 
    ra_2386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_945_inst_ack_0, ack => convolution3D_CP_1120_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	375 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	198 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_Update/$exit
      -- 
    ca_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_945_inst_ack_1, ack => convolution3D_CP_1120_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	185 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_Update/cr
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_update_start_
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_sample_completed_
      -- 
    ra_2400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_959_inst_ack_0, ack => convolution3D_CP_1120_elements(191)); -- 
    cr_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(191), ack => RPIPE_maxpool_input_pipe_959_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	196 
    -- CP-element group 192:  members (6) 
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_959_update_completed_
      -- 
    ca_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_959_inst_ack_1, ack => convolution3D_CP_1120_elements(192)); -- 
    rr_2427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(192), ack => type_cast_966_inst_req_0); -- 
    -- CP-element group 193:  join  transition  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_Sample/req
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_sample_start_
      -- 
    req_2413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(193), ack => WPIPE_maxpool_output_pipe_961_inst_req_0); -- 
    convolution3D_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(188) & convolution3D_CP_1120_elements(192);
      gj_convolution3D_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_update_start_
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_Update/req
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_sample_completed_
      -- 
    ack_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_961_inst_ack_0, ack => convolution3D_CP_1120_elements(194)); -- 
    req_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(194), ack => WPIPE_maxpool_output_pipe_961_inst_req_1); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	201 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_Update/ack
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/WPIPE_maxpool_output_pipe_961_update_completed_
      -- 
    ack_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_961_inst_ack_1, ack => convolution3D_CP_1120_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	192 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_Sample/ra
      -- 
    ra_2428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_966_inst_ack_0, ack => convolution3D_CP_1120_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	375 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_Update/ca
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_Update/$exit
      -- 
    ca_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_966_inst_ack_1, ack => convolution3D_CP_1120_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	142 
    -- CP-element group 198: 	148 
    -- CP-element group 198: 	155 
    -- CP-element group 198: 	162 
    -- CP-element group 198: 	169 
    -- CP-element group 198: 	176 
    -- CP-element group 198: 	183 
    -- CP-element group 198: 	190 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/word_access_start/word_0/rr
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/word_access_start/word_0/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/word_access_start/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/ptr_deref_974_Split/split_ack
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/ptr_deref_974_Split/split_req
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/ptr_deref_974_Split/$exit
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/ptr_deref_974_Split/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_sample_start_
      -- 
    rr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(198), ack => ptr_deref_974_store_0_req_0); -- 
    convolution3D_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(142) & convolution3D_CP_1120_elements(148) & convolution3D_CP_1120_elements(155) & convolution3D_CP_1120_elements(162) & convolution3D_CP_1120_elements(169) & convolution3D_CP_1120_elements(176) & convolution3D_CP_1120_elements(183) & convolution3D_CP_1120_elements(190) & convolution3D_CP_1120_elements(197);
      gj_convolution3D_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (5) 
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/word_access_start/word_0/ra
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/word_access_start/word_0/$exit
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/word_access_start/$exit
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_sample_completed_
      -- 
    ra_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_974_store_0_ack_0, ack => convolution3D_CP_1120_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	375 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (5) 
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Update/word_access_complete/word_0/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Update/word_access_complete/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Update/word_access_complete/word_0/ca
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_update_completed_
      -- 
    ca_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_974_store_0_ack_1, ack => convolution3D_CP_1120_elements(200)); -- 
    -- CP-element group 201:  branch  join  transition  place  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	139 
    -- CP-element group 201: 	195 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (10) 
      -- CP-element group 201: 	 branch_block_stmt_436/if_stmt_988_eval_test/$entry
      -- CP-element group 201: 	 branch_block_stmt_436/if_stmt_988_eval_test/$exit
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987__exit__
      -- CP-element group 201: 	 branch_block_stmt_436/if_stmt_988__entry__
      -- CP-element group 201: 	 branch_block_stmt_436/if_stmt_988_else_link/$entry
      -- CP-element group 201: 	 branch_block_stmt_436/if_stmt_988_dead_link/$entry
      -- CP-element group 201: 	 branch_block_stmt_436/R_exitcond32_989_place
      -- CP-element group 201: 	 branch_block_stmt_436/if_stmt_988_if_link/$entry
      -- CP-element group 201: 	 branch_block_stmt_436/if_stmt_988_eval_test/branch_req
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/$exit
      -- 
    branch_req_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(201), ack => if_stmt_988_branch_req_0); -- 
    convolution3D_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(139) & convolution3D_CP_1120_elements(195) & convolution3D_CP_1120_elements(200);
      gj_convolution3D_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	377 
    -- CP-element group 202: 	378 
    -- CP-element group 202:  members (24) 
      -- CP-element group 202: 	 branch_block_stmt_436/merge_stmt_994__exit__
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1016__entry__
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1016__exit__
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1016/$exit
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1016/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/if_stmt_988_if_link/if_choice_transition
      -- CP-element group 202: 	 branch_block_stmt_436/if_stmt_988_if_link/$exit
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 202: 	 branch_block_stmt_436/merge_stmt_994_PhiReqMerge
      -- CP-element group 202: 	 branch_block_stmt_436/merge_stmt_994_PhiAck/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/merge_stmt_994_PhiAck/$exit
      -- CP-element group 202: 	 branch_block_stmt_436/merge_stmt_994_PhiAck/dummy
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/Sample/rr
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_988_branch_ack_1, ack => convolution3D_CP_1120_elements(202)); -- 
    rr_3885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(202), ack => type_cast_1022_inst_req_0); -- 
    cr_3890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(202), ack => type_cast_1022_inst_req_1); -- 
    -- CP-element group 203:  fork  transition  place  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	371 
    -- CP-element group 203: 	372 
    -- CP-element group 203:  members (12) 
      -- CP-element group 203: 	 branch_block_stmt_436/if_stmt_988_else_link/else_choice_transition
      -- CP-element group 203: 	 branch_block_stmt_436/if_stmt_988_else_link/$exit
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/Sample/rr
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_988_branch_ack_0, ack => convolution3D_CP_1120_elements(203)); -- 
    rr_3831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(203), ack => type_cast_807_inst_req_0); -- 
    cr_3836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(203), ack => type_cast_807_inst_req_1); -- 
    -- CP-element group 204:  transition  place  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	381 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	400 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_436/if_stmt_1039_if_link/if_choice_transition
      -- CP-element group 204: 	 branch_block_stmt_436/if_stmt_1039_if_link/$exit
      -- CP-element group 204: 	 branch_block_stmt_436/forx_xend_ifx_xend
      -- CP-element group 204: 	 branch_block_stmt_436/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 204: 	 branch_block_stmt_436/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1039_branch_ack_1, ack => convolution3D_CP_1120_elements(204)); -- 
    -- CP-element group 205:  merge  fork  transition  place  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	381 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	382 
    -- CP-element group 205: 	383 
    -- CP-element group 205:  members (20) 
      -- CP-element group 205: 	 branch_block_stmt_436/merge_stmt_1045__exit__
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1057__entry__
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1057__exit__
      -- CP-element group 205: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1057/$exit
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1051_to_assign_stmt_1057/$entry
      -- CP-element group 205: 	 branch_block_stmt_436/if_stmt_1039_else_link/else_choice_transition
      -- CP-element group 205: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi
      -- CP-element group 205: 	 branch_block_stmt_436/if_stmt_1039_else_link/$exit
      -- CP-element group 205: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 205: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 205: 	 branch_block_stmt_436/merge_stmt_1045_PhiReqMerge
      -- CP-element group 205: 	 branch_block_stmt_436/merge_stmt_1045_PhiAck/$entry
      -- CP-element group 205: 	 branch_block_stmt_436/merge_stmt_1045_PhiAck/$exit
      -- CP-element group 205: 	 branch_block_stmt_436/merge_stmt_1045_PhiAck/dummy
      -- CP-element group 205: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 205: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/$entry
      -- CP-element group 205: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/$entry
      -- CP-element group 205: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/$entry
      -- CP-element group 205: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/$entry
      -- 
    else_choice_transition_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1039_branch_ack_0, ack => convolution3D_CP_1120_elements(205)); -- 
    -- CP-element group 206:  transition  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	395 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (6) 
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_Update/cr
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_Sample/ra
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_update_start_
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_sample_completed_
      -- 
    ra_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1088_inst_ack_0, ack => convolution3D_CP_1120_elements(206)); -- 
    cr_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(206), ack => RPIPE_maxpool_input_pipe_1088_inst_req_1); -- 
    -- CP-element group 207:  fork  transition  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207: 	210 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_Update/ca
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_Sample/req
      -- 
    ca_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1088_inst_ack_1, ack => convolution3D_CP_1120_elements(207)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(207), ack => WPIPE_maxpool_output_pipe_1090_inst_req_0); -- 
    rr_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(207), ack => type_cast_1095_inst_req_0); -- 
    -- CP-element group 208:  transition  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_update_start_
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_Update/req
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_Sample/ack
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1090_inst_ack_0, ack => convolution3D_CP_1120_elements(208)); -- 
    req_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(208), ack => WPIPE_maxpool_output_pipe_1090_inst_req_1); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	214 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_Update/ack
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/WPIPE_maxpool_output_pipe_1090_Update/$exit
      -- 
    ack_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1090_inst_ack_1, ack => convolution3D_CP_1120_elements(209)); -- 
    -- CP-element group 210:  transition  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	207 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_Sample/ra
      -- CP-element group 210: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_Sample/$exit
      -- CP-element group 210: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_sample_completed_
      -- 
    ra_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1095_inst_ack_0, ack => convolution3D_CP_1120_elements(210)); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	395 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	214 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_Update/ca
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_Update/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_update_completed_
      -- 
    ca_2575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1095_inst_ack_1, ack => convolution3D_CP_1120_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	395 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_Sample/ra
      -- CP-element group 212: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_Sample/$exit
      -- 
    ra_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_0, ack => convolution3D_CP_1120_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	395 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_Update/ca
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_Update/$exit
      -- 
    ca_2589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_1, ack => convolution3D_CP_1120_elements(213)); -- 
    -- CP-element group 214:  branch  join  transition  place  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	209 
    -- CP-element group 214: 	211 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (10) 
      -- CP-element group 214: 	 branch_block_stmt_436/R_cmpx_xi_1118_place
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116__exit__
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1117__entry__
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1117_else_link/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1117_if_link/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1117_eval_test/branch_req
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/$exit
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1117_eval_test/$exit
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1117_eval_test/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1117_dead_link/$entry
      -- 
    branch_req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(214), ack => if_stmt_1117_branch_req_0); -- 
    convolution3D_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(209) & convolution3D_CP_1120_elements(211) & convolution3D_CP_1120_elements(213);
      gj_convolution3D_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  fork  transition  place  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	385 
    -- CP-element group 215: 	386 
    -- CP-element group 215: 	388 
    -- CP-element group 215: 	389 
    -- CP-element group 215:  members (20) 
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 215: 	 branch_block_stmt_436/if_stmt_1117_if_link/if_choice_transition
      -- CP-element group 215: 	 branch_block_stmt_436/if_stmt_1117_if_link/$exit
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/Sample/rr
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/Update/cr
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/Sample/rr
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1117_branch_ack_1, ack => convolution3D_CP_1120_elements(215)); -- 
    rr_3947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(215), ack => type_cast_1066_inst_req_0); -- 
    cr_3952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(215), ack => type_cast_1066_inst_req_1); -- 
    rr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(215), ack => type_cast_1073_inst_req_0); -- 
    cr_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(215), ack => type_cast_1073_inst_req_1); -- 
    -- CP-element group 216:  fork  transition  place  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	396 
    -- CP-element group 216: 	397 
    -- CP-element group 216:  members (12) 
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 216: 	 branch_block_stmt_436/if_stmt_1117_else_link/else_choice_transition
      -- CP-element group 216: 	 branch_block_stmt_436/if_stmt_1117_else_link/$exit
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/Sample/rr
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1117_branch_ack_0, ack => convolution3D_CP_1120_elements(216)); -- 
    rr_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(216), ack => type_cast_1127_inst_req_0); -- 
    cr_4011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(216), ack => type_cast_1127_inst_req_1); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	399 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	223 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_sample_complete
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_Sample/ack
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_Sample/$exit
      -- 
    ack_2637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1156_index_offset_ack_0, ack => convolution3D_CP_1120_elements(217)); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	399 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (11) 
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_root_address_calculated
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_offset_calculated
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_request/req
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_Update/ack
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_request/$entry
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_base_plus_offset/sum_rename_ack
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_base_plus_offset/sum_rename_req
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_base_plus_offset/$exit
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_base_plus_offset/$entry
      -- 
    ack_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1156_index_offset_ack_1, ack => convolution3D_CP_1120_elements(218)); -- 
    req_2651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => addr_of_1157_final_reg_req_0); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_request/ack
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_request/$exit
      -- 
    ack_2652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1157_final_reg_ack_0, ack => convolution3D_CP_1120_elements(219)); -- 
    -- CP-element group 220:  join  fork  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	399 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (28) 
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_addr_resize/$exit
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_addr_resize/base_resize_req
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_addr_resize/base_resize_ack
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_plus_offset/$entry
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_addr_resize/$entry
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_address_resized
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_root_address_calculated
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_word_address_calculated
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_address_calculated
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/word_access_start/word_0/rr
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_complete/ack
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_complete/$exit
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/word_access_start/word_0/$entry
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/word_access_start/$entry
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/ptr_deref_1160_Split/split_ack
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/ptr_deref_1160_Split/split_req
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/ptr_deref_1160_Split/$exit
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/ptr_deref_1160_Split/$entry
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_word_addrgen/root_register_ack
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_word_addrgen/root_register_req
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_word_addrgen/$exit
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_word_addrgen/$entry
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_plus_offset/sum_rename_ack
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_plus_offset/sum_rename_req
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_base_plus_offset/$exit
      -- 
    ack_2657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1157_final_reg_ack_1, ack => convolution3D_CP_1120_elements(220)); -- 
    rr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(220), ack => ptr_deref_1160_store_0_req_0); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (5) 
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/word_access_start/word_0/ra
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/word_access_start/word_0/$exit
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/word_access_start/$exit
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Sample/$exit
      -- 
    ra_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1160_store_0_ack_0, ack => convolution3D_CP_1120_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	399 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (5) 
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Update/word_access_complete/word_0/ca
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Update/word_access_complete/word_0/$exit
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Update/word_access_complete/$exit
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_update_completed_
      -- 
    ca_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1160_store_0_ack_1, ack => convolution3D_CP_1120_elements(222)); -- 
    -- CP-element group 223:  join  transition  place  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	217 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	400 
    -- CP-element group 223:  members (5) 
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/$exit
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162__exit__
      -- CP-element group 223: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 223: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 223: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(217) & convolution3D_CP_1120_elements(222);
      gj_convolution3D_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	400 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_Sample/ra
      -- CP-element group 224: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_Sample/$exit
      -- 
    ra_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_0, ack => convolution3D_CP_1120_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	400 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	232 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_Update/ca
      -- CP-element group 225: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_update_completed_
      -- 
    ca_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_1, ack => convolution3D_CP_1120_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	400 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_Sample/ra
      -- 
    ra_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_0, ack => convolution3D_CP_1120_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	400 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	232 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_Update/ca
      -- 
    ca_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_1, ack => convolution3D_CP_1120_elements(227)); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	400 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_Sample/ra
      -- 
    ra_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1175_inst_ack_0, ack => convolution3D_CP_1120_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	400 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	232 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_Update/ca
      -- 
    ca_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1175_inst_ack_1, ack => convolution3D_CP_1120_elements(229)); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	400 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_Sample/ra
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1179_inst_ack_0, ack => convolution3D_CP_1120_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	400 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_Update/ca
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1179_inst_ack_1, ack => convolution3D_CP_1120_elements(231)); -- 
    -- CP-element group 232:  branch  join  transition  place  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	225 
    -- CP-element group 232: 	227 
    -- CP-element group 232: 	229 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (10) 
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/$exit
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216__exit__
      -- CP-element group 232: 	 branch_block_stmt_436/if_stmt_1217__entry__
      -- CP-element group 232: 	 branch_block_stmt_436/if_stmt_1217_dead_link/$entry
      -- CP-element group 232: 	 branch_block_stmt_436/if_stmt_1217_eval_test/$entry
      -- CP-element group 232: 	 branch_block_stmt_436/if_stmt_1217_eval_test/$exit
      -- CP-element group 232: 	 branch_block_stmt_436/if_stmt_1217_eval_test/branch_req
      -- CP-element group 232: 	 branch_block_stmt_436/R_cmp255443_1218_place
      -- CP-element group 232: 	 branch_block_stmt_436/if_stmt_1217_if_link/$entry
      -- CP-element group 232: 	 branch_block_stmt_436/if_stmt_1217_else_link/$entry
      -- 
    branch_req_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(232), ack => if_stmt_1217_branch_req_0); -- 
    convolution3D_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(225) & convolution3D_CP_1120_elements(227) & convolution3D_CP_1120_elements(229) & convolution3D_CP_1120_elements(231);
      gj_convolution3D_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: 	236 
    -- CP-element group 233: 	237 
    -- CP-element group 233: 	238 
    -- CP-element group 233: 	239 
    -- CP-element group 233: 	240 
    -- CP-element group 233: 	241 
    -- CP-element group 233: 	242 
    -- CP-element group 233: 	245 
    -- CP-element group 233: 	247 
    -- CP-element group 233:  members (42) 
      -- CP-element group 233: 	 branch_block_stmt_436/merge_stmt_1223__exit__
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294__entry__
      -- CP-element group 233: 	 branch_block_stmt_436/if_stmt_1217_if_link/$exit
      -- CP-element group 233: 	 branch_block_stmt_436/if_stmt_1217_if_link/if_choice_transition
      -- CP-element group 233: 	 branch_block_stmt_436/ifx_xend_bbx_xnph
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_update_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_Sample/rr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_update_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_Sample/rr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_update_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_Sample/rr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_update_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_Sample/rr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_update_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_update_start_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_436/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 233: 	 branch_block_stmt_436/merge_stmt_1223_PhiReqMerge
      -- CP-element group 233: 	 branch_block_stmt_436/merge_stmt_1223_PhiAck/$entry
      -- CP-element group 233: 	 branch_block_stmt_436/merge_stmt_1223_PhiAck/$exit
      -- CP-element group 233: 	 branch_block_stmt_436/merge_stmt_1223_PhiAck/dummy
      -- 
    if_choice_transition_2779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1217_branch_ack_1, ack => convolution3D_CP_1120_elements(233)); -- 
    rr_2796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1238_inst_req_0); -- 
    cr_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1238_inst_req_1); -- 
    rr_2810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1242_inst_req_0); -- 
    cr_2815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1242_inst_req_1); -- 
    rr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1251_inst_req_0); -- 
    cr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1251_inst_req_1); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1260_inst_req_0); -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1260_inst_req_1); -- 
    cr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1269_inst_req_1); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(233), ack => type_cast_1274_inst_req_1); -- 
    -- CP-element group 234:  transition  place  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	410 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_436/if_stmt_1217_else_link/$exit
      -- CP-element group 234: 	 branch_block_stmt_436/if_stmt_1217_else_link/else_choice_transition
      -- CP-element group 234: 	 branch_block_stmt_436/ifx_xend_forx_xend341
      -- CP-element group 234: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1515/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$entry
      -- 
    else_choice_transition_2783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1217_branch_ack_0, ack => convolution3D_CP_1120_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_Sample/ra
      -- 
    ra_2797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => convolution3D_CP_1120_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	233 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	243 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1238_Update/ca
      -- 
    ca_2802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => convolution3D_CP_1120_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	233 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_Sample/ra
      -- 
    ra_2811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1242_inst_ack_0, ack => convolution3D_CP_1120_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	233 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	243 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1242_Update/ca
      -- 
    ca_2816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1242_inst_ack_1, ack => convolution3D_CP_1120_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	233 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_Sample/ra
      -- 
    ra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_0, ack => convolution3D_CP_1120_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	233 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	243 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1251_Update/ca
      -- 
    ca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_1, ack => convolution3D_CP_1120_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	233 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_Sample/ra
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1260_inst_ack_0, ack => convolution3D_CP_1120_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	233 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1260_Update/ca
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1260_inst_ack_1, ack => convolution3D_CP_1120_elements(242)); -- 
    -- CP-element group 243:  join  transition  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	236 
    -- CP-element group 243: 	238 
    -- CP-element group 243: 	240 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_Sample/rr
      -- 
    rr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(243), ack => type_cast_1269_inst_req_0); -- 
    convolution3D_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(236) & convolution3D_CP_1120_elements(238) & convolution3D_CP_1120_elements(240) & convolution3D_CP_1120_elements(242);
      gj_convolution3D_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_Sample/ra
      -- 
    ra_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_0, ack => convolution3D_CP_1120_elements(244)); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	233 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1269_Update/ca
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_Sample/rr
      -- 
    ca_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_1, ack => convolution3D_CP_1120_elements(245)); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(245), ack => type_cast_1274_inst_req_0); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_Sample/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1274_inst_ack_0, ack => convolution3D_CP_1120_elements(246)); -- 
    -- CP-element group 247:  transition  place  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	233 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	401 
    -- CP-element group 247:  members (9) 
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294__exit__
      -- CP-element group 247: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/$exit
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1294/type_cast_1274_Update/ca
      -- CP-element group 247: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/$entry
      -- CP-element group 247: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1297/$entry
      -- CP-element group 247: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/$entry
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1274_inst_ack_1, ack => convolution3D_CP_1120_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	406 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	310 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_sample_complete
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_Sample/ack
      -- 
    ack_2901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1309_index_offset_ack_0, ack => convolution3D_CP_1120_elements(248)); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	406 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (11) 
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_root_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_offset_calculated
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_Update/ack
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_base_plus_offset/$entry
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_base_plus_offset/$exit
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_base_plus_offset/sum_rename_req
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_base_plus_offset/sum_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_request/$entry
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_request/req
      -- 
    ack_2906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1309_index_offset_ack_1, ack => convolution3D_CP_1120_elements(249)); -- 
    req_2915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => addr_of_1310_final_reg_req_0); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_request/$exit
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_request/ack
      -- 
    ack_2916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1310_final_reg_ack_0, ack => convolution3D_CP_1120_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	406 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	307 
    -- CP-element group 251:  members (19) 
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_complete/$exit
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_complete/ack
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_address_calculated
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_word_address_calculated
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_root_address_calculated
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_address_resized
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_addr_resize/$entry
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_addr_resize/$exit
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_addr_resize/base_resize_req
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_addr_resize/base_resize_ack
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_plus_offset/$entry
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_plus_offset/$exit
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_plus_offset/sum_rename_req
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_base_plus_offset/sum_rename_ack
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_word_addrgen/$entry
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_word_addrgen/$exit
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_word_addrgen/root_register_req
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_word_addrgen/root_register_ack
      -- 
    ack_2921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1310_final_reg_ack_1, ack => convolution3D_CP_1120_elements(251)); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	406 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_update_start_
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_Sample/ra
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_Update/$entry
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_Update/cr
      -- 
    ra_2930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1313_inst_ack_0, ack => convolution3D_CP_1120_elements(252)); -- 
    cr_2934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(252), ack => RPIPE_maxpool_input_pipe_1313_inst_req_1); -- 
    -- CP-element group 253:  fork  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253: 	256 
    -- CP-element group 253: 	258 
    -- CP-element group 253:  members (12) 
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_Update/ca
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_Sample/req
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_Sample/rr
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_Sample/rr
      -- 
    ca_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1313_inst_ack_1, ack => convolution3D_CP_1120_elements(253)); -- 
    req_2943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(253), ack => WPIPE_maxpool_output_pipe_1315_inst_req_0); -- 
    rr_2957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(253), ack => type_cast_1320_inst_req_0); -- 
    rr_2971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(253), ack => RPIPE_maxpool_input_pipe_1329_inst_req_0); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_update_start_
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_Sample/ack
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_Update/req
      -- 
    ack_2944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1315_inst_ack_0, ack => convolution3D_CP_1120_elements(254)); -- 
    req_2948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(254), ack => WPIPE_maxpool_output_pipe_1315_inst_req_1); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	260 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1315_Update/ack
      -- 
    ack_2949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1315_inst_ack_1, ack => convolution3D_CP_1120_elements(255)); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	253 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_Sample/ra
      -- 
    ra_2958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_0, ack => convolution3D_CP_1120_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	406 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	307 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_Update/ca
      -- 
    ca_2963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_1, ack => convolution3D_CP_1120_elements(257)); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	253 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_sample_completed_
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_update_start_
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_Sample/ra
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_Update/cr
      -- 
    ra_2972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1329_inst_ack_0, ack => convolution3D_CP_1120_elements(258)); -- 
    cr_2976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(258), ack => RPIPE_maxpool_input_pipe_1329_inst_req_1); -- 
    -- CP-element group 259:  fork  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259: 	263 
    -- CP-element group 259: 	265 
    -- CP-element group 259:  members (9) 
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1329_Update/ca
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_Sample/rr
      -- 
    ca_2977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1329_inst_ack_1, ack => convolution3D_CP_1120_elements(259)); -- 
    rr_2999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(259), ack => type_cast_1336_inst_req_0); -- 
    rr_3013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(259), ack => RPIPE_maxpool_input_pipe_1350_inst_req_0); -- 
    -- CP-element group 260:  join  transition  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	255 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_Sample/req
      -- 
    req_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(260), ack => WPIPE_maxpool_output_pipe_1331_inst_req_0); -- 
    convolution3D_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(255) & convolution3D_CP_1120_elements(259);
      gj_convolution3D_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_update_start_
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_Update/req
      -- 
    ack_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1331_inst_ack_0, ack => convolution3D_CP_1120_elements(261)); -- 
    req_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(261), ack => WPIPE_maxpool_output_pipe_1331_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	267 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1331_Update/ack
      -- 
    ack_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1331_inst_ack_1, ack => convolution3D_CP_1120_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	259 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_Sample/ra
      -- 
    ra_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1336_inst_ack_0, ack => convolution3D_CP_1120_elements(263)); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	406 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	307 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_Update/ca
      -- 
    ca_3005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1336_inst_ack_1, ack => convolution3D_CP_1120_elements(264)); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	259 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_update_start_
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_Sample/ra
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_Update/cr
      -- 
    ra_3014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1350_inst_ack_0, ack => convolution3D_CP_1120_elements(265)); -- 
    cr_3018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(265), ack => RPIPE_maxpool_input_pipe_1350_inst_req_1); -- 
    -- CP-element group 266:  fork  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266: 	270 
    -- CP-element group 266: 	272 
    -- CP-element group 266:  members (9) 
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1350_Update/ca
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_Sample/rr
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_Sample/rr
      -- 
    ca_3019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1350_inst_ack_1, ack => convolution3D_CP_1120_elements(266)); -- 
    rr_3041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(266), ack => type_cast_1357_inst_req_0); -- 
    rr_3055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(266), ack => RPIPE_maxpool_input_pipe_1371_inst_req_0); -- 
    -- CP-element group 267:  join  transition  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	262 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_Sample/req
      -- 
    req_3027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(267), ack => WPIPE_maxpool_output_pipe_1352_inst_req_0); -- 
    convolution3D_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(262) & convolution3D_CP_1120_elements(266);
      gj_convolution3D_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_update_start_
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_Sample/ack
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_Update/req
      -- 
    ack_3028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1352_inst_ack_0, ack => convolution3D_CP_1120_elements(268)); -- 
    req_3032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(268), ack => WPIPE_maxpool_output_pipe_1352_inst_req_1); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	274 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1352_Update/ack
      -- 
    ack_3033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1352_inst_ack_1, ack => convolution3D_CP_1120_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	266 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_Sample/ra
      -- 
    ra_3042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1357_inst_ack_0, ack => convolution3D_CP_1120_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	406 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	307 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_Update/ca
      -- 
    ca_3047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1357_inst_ack_1, ack => convolution3D_CP_1120_elements(271)); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	266 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_update_start_
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_Sample/ra
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_Update/cr
      -- 
    ra_3056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1371_inst_ack_0, ack => convolution3D_CP_1120_elements(272)); -- 
    cr_3060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(272), ack => RPIPE_maxpool_input_pipe_1371_inst_req_1); -- 
    -- CP-element group 273:  fork  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273: 	277 
    -- CP-element group 273: 	279 
    -- CP-element group 273:  members (9) 
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1371_Update/ca
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_sample_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_Sample/rr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_sample_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_Sample/rr
      -- 
    ca_3061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1371_inst_ack_1, ack => convolution3D_CP_1120_elements(273)); -- 
    rr_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_1378_inst_req_0); -- 
    rr_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => RPIPE_maxpool_input_pipe_1392_inst_req_0); -- 
    -- CP-element group 274:  join  transition  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	269 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_Sample/req
      -- 
    req_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(274), ack => WPIPE_maxpool_output_pipe_1373_inst_req_0); -- 
    convolution3D_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(269) & convolution3D_CP_1120_elements(273);
      gj_convolution3D_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_sample_completed_
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_update_start_
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_Update/req
      -- 
    ack_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1373_inst_ack_0, ack => convolution3D_CP_1120_elements(275)); -- 
    req_3074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(275), ack => WPIPE_maxpool_output_pipe_1373_inst_req_1); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	281 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1373_Update/ack
      -- 
    ack_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1373_inst_ack_1, ack => convolution3D_CP_1120_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	273 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_Sample/ra
      -- 
    ra_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_0, ack => convolution3D_CP_1120_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	406 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	307 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_Update/ca
      -- 
    ca_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_1, ack => convolution3D_CP_1120_elements(278)); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	273 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_update_start_
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_Update/cr
      -- 
    ra_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1392_inst_ack_0, ack => convolution3D_CP_1120_elements(279)); -- 
    cr_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(279), ack => RPIPE_maxpool_input_pipe_1392_inst_req_1); -- 
    -- CP-element group 280:  fork  transition  input  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280: 	284 
    -- CP-element group 280: 	286 
    -- CP-element group 280:  members (9) 
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1392_Update/ca
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_Sample/rr
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_Sample/rr
      -- 
    ca_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1392_inst_ack_1, ack => convolution3D_CP_1120_elements(280)); -- 
    rr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(280), ack => type_cast_1399_inst_req_0); -- 
    rr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(280), ack => RPIPE_maxpool_input_pipe_1413_inst_req_0); -- 
    -- CP-element group 281:  join  transition  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	276 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_Sample/req
      -- 
    req_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(281), ack => WPIPE_maxpool_output_pipe_1394_inst_req_0); -- 
    convolution3D_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(276) & convolution3D_CP_1120_elements(280);
      gj_convolution3D_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (6) 
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_sample_completed_
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_update_start_
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_Sample/ack
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_Update/$entry
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_Update/req
      -- 
    ack_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1394_inst_ack_0, ack => convolution3D_CP_1120_elements(282)); -- 
    req_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(282), ack => WPIPE_maxpool_output_pipe_1394_inst_req_1); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	288 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_update_completed_
      -- CP-element group 283: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1394_Update/ack
      -- 
    ack_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1394_inst_ack_1, ack => convolution3D_CP_1120_elements(283)); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	280 
    -- CP-element group 284: successors 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_Sample/ra
      -- 
    ra_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1399_inst_ack_0, ack => convolution3D_CP_1120_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	406 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	307 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_Update/ca
      -- 
    ca_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1399_inst_ack_1, ack => convolution3D_CP_1120_elements(285)); -- 
    -- CP-element group 286:  transition  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	280 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (6) 
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_update_start_
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_Update/$entry
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_Update/cr
      -- 
    ra_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1413_inst_ack_0, ack => convolution3D_CP_1120_elements(286)); -- 
    cr_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(286), ack => RPIPE_maxpool_input_pipe_1413_inst_req_1); -- 
    -- CP-element group 287:  fork  transition  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	293 
    -- CP-element group 287: 	288 
    -- CP-element group 287: 	291 
    -- CP-element group 287:  members (9) 
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1413_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_Sample/rr
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_Sample/rr
      -- 
    ca_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1413_inst_ack_1, ack => convolution3D_CP_1120_elements(287)); -- 
    rr_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(287), ack => RPIPE_maxpool_input_pipe_1434_inst_req_0); -- 
    rr_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(287), ack => type_cast_1420_inst_req_0); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	283 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_Sample/req
      -- 
    req_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(288), ack => WPIPE_maxpool_output_pipe_1415_inst_req_0); -- 
    convolution3D_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(283) & convolution3D_CP_1120_elements(287);
      gj_convolution3D_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_sample_completed_
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_update_start_
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_Update/req
      -- 
    ack_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1415_inst_ack_0, ack => convolution3D_CP_1120_elements(289)); -- 
    req_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(289), ack => WPIPE_maxpool_output_pipe_1415_inst_req_1); -- 
    -- CP-element group 290:  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	295 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1415_Update/ack
      -- 
    ack_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1415_inst_ack_1, ack => convolution3D_CP_1120_elements(290)); -- 
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	287 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_Sample/ra
      -- 
    ra_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1420_inst_ack_0, ack => convolution3D_CP_1120_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	406 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	307 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_Update/ca
      -- 
    ca_3173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1420_inst_ack_1, ack => convolution3D_CP_1120_elements(292)); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	287 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_update_start_
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_Sample/ra
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_Update/cr
      -- 
    ra_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1434_inst_ack_0, ack => convolution3D_CP_1120_elements(293)); -- 
    cr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(293), ack => RPIPE_maxpool_input_pipe_1434_inst_req_1); -- 
    -- CP-element group 294:  fork  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294: 	298 
    -- CP-element group 294: 	300 
    -- CP-element group 294:  members (9) 
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1434_Update/ca
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_Sample/rr
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_Sample/rr
      -- 
    ca_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1434_inst_ack_1, ack => convolution3D_CP_1120_elements(294)); -- 
    rr_3209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(294), ack => type_cast_1441_inst_req_0); -- 
    rr_3223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(294), ack => RPIPE_maxpool_input_pipe_1455_inst_req_0); -- 
    -- CP-element group 295:  join  transition  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: 	290 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_Sample/req
      -- 
    req_3195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(295), ack => WPIPE_maxpool_output_pipe_1436_inst_req_0); -- 
    convolution3D_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(294) & convolution3D_CP_1120_elements(290);
      gj_convolution3D_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  transition  input  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (6) 
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_sample_completed_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_update_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_Sample/ack
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_Update/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_Update/req
      -- 
    ack_3196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1436_inst_ack_0, ack => convolution3D_CP_1120_elements(296)); -- 
    req_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => WPIPE_maxpool_output_pipe_1436_inst_req_1); -- 
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	302 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_update_completed_
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1436_Update/ack
      -- 
    ack_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1436_inst_ack_1, ack => convolution3D_CP_1120_elements(297)); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	294 
    -- CP-element group 298: successors 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_sample_completed_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_Sample/$exit
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_Sample/ra
      -- 
    ra_3210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1441_inst_ack_0, ack => convolution3D_CP_1120_elements(298)); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	406 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	307 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_update_completed_
      -- CP-element group 299: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_Update/$exit
      -- CP-element group 299: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_Update/ca
      -- 
    ca_3215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1441_inst_ack_1, ack => convolution3D_CP_1120_elements(299)); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	294 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_update_start_
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_Sample/ra
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_Update/cr
      -- 
    ra_3224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1455_inst_ack_0, ack => convolution3D_CP_1120_elements(300)); -- 
    cr_3228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(300), ack => RPIPE_maxpool_input_pipe_1455_inst_req_1); -- 
    -- CP-element group 301:  fork  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	305 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1455_Update/ca
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_Sample/rr
      -- 
    ca_3229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1455_inst_ack_1, ack => convolution3D_CP_1120_elements(301)); -- 
    rr_3251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(301), ack => type_cast_1462_inst_req_0); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	297 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_Sample/req
      -- 
    req_3237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => WPIPE_maxpool_output_pipe_1457_inst_req_0); -- 
    convolution3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(297) & convolution3D_CP_1120_elements(301);
      gj_convolution3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_update_start_
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_Update/req
      -- 
    ack_3238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1457_inst_ack_0, ack => convolution3D_CP_1120_elements(303)); -- 
    req_3242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(303), ack => WPIPE_maxpool_output_pipe_1457_inst_req_1); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	310 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/WPIPE_maxpool_output_pipe_1457_Update/ack
      -- 
    ack_3243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1457_inst_ack_1, ack => convolution3D_CP_1120_elements(304)); -- 
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	301 
    -- CP-element group 305: successors 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_Sample/ra
      -- 
    ra_3252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1462_inst_ack_0, ack => convolution3D_CP_1120_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	406 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_Update/ca
      -- 
    ca_3257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1462_inst_ack_1, ack => convolution3D_CP_1120_elements(306)); -- 
    -- CP-element group 307:  join  transition  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	292 
    -- CP-element group 307: 	306 
    -- CP-element group 307: 	299 
    -- CP-element group 307: 	251 
    -- CP-element group 307: 	257 
    -- CP-element group 307: 	264 
    -- CP-element group 307: 	271 
    -- CP-element group 307: 	278 
    -- CP-element group 307: 	285 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (9) 
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/word_access_start/word_0/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/word_access_start/word_0/rr
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/word_access_start/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/ptr_deref_1470_Split/split_ack
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/ptr_deref_1470_Split/split_req
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/ptr_deref_1470_Split/$exit
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/ptr_deref_1470_Split/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_sample_start_
      -- CP-element group 307: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/$entry
      -- 
    rr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(307), ack => ptr_deref_1470_store_0_req_0); -- 
    convolution3D_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(292) & convolution3D_CP_1120_elements(306) & convolution3D_CP_1120_elements(299) & convolution3D_CP_1120_elements(251) & convolution3D_CP_1120_elements(257) & convolution3D_CP_1120_elements(264) & convolution3D_CP_1120_elements(271) & convolution3D_CP_1120_elements(278) & convolution3D_CP_1120_elements(285);
      gj_convolution3D_cp_element_group_307 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308:  members (5) 
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/word_access_start/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/word_access_start/word_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/word_access_start/word_0/ra
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_sample_completed_
      -- CP-element group 308: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Sample/$exit
      -- 
    ra_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1470_store_0_ack_0, ack => convolution3D_CP_1120_elements(308)); -- 
    -- CP-element group 309:  transition  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	406 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (5) 
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Update/$exit
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Update/word_access_complete/word_0/ca
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Update/word_access_complete/word_0/$exit
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Update/word_access_complete/$exit
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_update_completed_
      -- 
    ca_3307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1470_store_0_ack_1, ack => convolution3D_CP_1120_elements(309)); -- 
    -- CP-element group 310:  branch  join  transition  place  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: 	304 
    -- CP-element group 310: 	248 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (10) 
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483__exit__
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1484__entry__
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1484_if_link/$entry
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1484_else_link/$entry
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1484_eval_test/branch_req
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1484_eval_test/$exit
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1484_eval_test/$entry
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1484_dead_link/$entry
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/$exit
      -- CP-element group 310: 	 branch_block_stmt_436/R_exitcond_1485_place
      -- 
    branch_req_3315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(310), ack => if_stmt_1484_branch_req_0); -- 
    convolution3D_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(309) & convolution3D_CP_1120_elements(304) & convolution3D_CP_1120_elements(248);
      gj_convolution3D_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	407 
    -- CP-element group 311: 	408 
    -- CP-element group 311:  members (24) 
      -- CP-element group 311: 	 branch_block_stmt_436/merge_stmt_1490__exit__
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1497_to_assign_stmt_1512__entry__
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1497_to_assign_stmt_1512__exit__
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341
      -- CP-element group 311: 	 branch_block_stmt_436/if_stmt_1484_if_link/$exit
      -- CP-element group 311: 	 branch_block_stmt_436/if_stmt_1484_if_link/if_choice_transition
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xbody257_forx_xcond250x_xforx_xend341_crit_edge
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1497_to_assign_stmt_1512/$exit
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1497_to_assign_stmt_1512/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xbody257_forx_xcond250x_xforx_xend341_crit_edge_PhiReq/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xbody257_forx_xcond250x_xforx_xend341_crit_edge_PhiReq/$exit
      -- CP-element group 311: 	 branch_block_stmt_436/merge_stmt_1490_PhiReqMerge
      -- CP-element group 311: 	 branch_block_stmt_436/merge_stmt_1490_PhiAck/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/merge_stmt_1490_PhiAck/$exit
      -- CP-element group 311: 	 branch_block_stmt_436/merge_stmt_1490_PhiAck/dummy
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/rr
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1484_branch_ack_1, ack => convolution3D_CP_1120_elements(311)); -- 
    rr_4114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(311), ack => type_cast_1521_inst_req_0); -- 
    cr_4119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(311), ack => type_cast_1521_inst_req_1); -- 
    -- CP-element group 312:  fork  transition  place  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	402 
    -- CP-element group 312: 	403 
    -- CP-element group 312:  members (12) 
      -- CP-element group 312: 	 branch_block_stmt_436/if_stmt_1484_else_link/$exit
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257
      -- CP-element group 312: 	 branch_block_stmt_436/if_stmt_1484_else_link/else_choice_transition
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/$entry
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/$entry
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/$entry
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/$entry
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/$entry
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Sample/rr
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1484_branch_ack_0, ack => convolution3D_CP_1120_elements(312)); -- 
    rr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(312), ack => type_cast_1303_inst_req_0); -- 
    cr_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(312), ack => type_cast_1303_inst_req_1); -- 
    -- CP-element group 313:  transition  place  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	412 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	431 
    -- CP-element group 313:  members (5) 
      -- CP-element group 313: 	 branch_block_stmt_436/forx_xend341_ifx_xend353
      -- CP-element group 313: 	 branch_block_stmt_436/if_stmt_1535_if_link/if_choice_transition
      -- CP-element group 313: 	 branch_block_stmt_436/if_stmt_1535_if_link/$exit
      -- CP-element group 313: 	 branch_block_stmt_436/forx_xend341_ifx_xend353_PhiReq/$entry
      -- CP-element group 313: 	 branch_block_stmt_436/forx_xend341_ifx_xend353_PhiReq/$exit
      -- 
    if_choice_transition_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1535_branch_ack_1, ack => convolution3D_CP_1120_elements(313)); -- 
    -- CP-element group 314:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	412 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (18) 
      -- CP-element group 314: 	 branch_block_stmt_436/merge_stmt_1541__exit__
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557__entry__
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_Sample/rr
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_update_start_
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_Sample/$entry
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xend341_bbx_xnphx_xi420
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_sample_start_
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/$entry
      -- CP-element group 314: 	 branch_block_stmt_436/if_stmt_1535_else_link/else_choice_transition
      -- CP-element group 314: 	 branch_block_stmt_436/if_stmt_1535_else_link/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_Update/cr
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_Update/$entry
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xend341_bbx_xnphx_xi420_PhiReq/$entry
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xend341_bbx_xnphx_xi420_PhiReq/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/merge_stmt_1541_PhiReqMerge
      -- CP-element group 314: 	 branch_block_stmt_436/merge_stmt_1541_PhiAck/$entry
      -- CP-element group 314: 	 branch_block_stmt_436/merge_stmt_1541_PhiAck/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/merge_stmt_1541_PhiAck/dummy
      -- 
    else_choice_transition_3349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1535_branch_ack_0, ack => convolution3D_CP_1120_elements(314)); -- 
    rr_3362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(314), ack => type_cast_1550_inst_req_0); -- 
    cr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(314), ack => type_cast_1550_inst_req_1); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_Sample/ra
      -- 
    ra_3363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1550_inst_ack_0, ack => convolution3D_CP_1120_elements(315)); -- 
    -- CP-element group 316:  fork  transition  place  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	414 
    -- CP-element group 316: 	413 
    -- CP-element group 316:  members (11) 
      -- CP-element group 316: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557__exit__
      -- CP-element group 316: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429
      -- CP-element group 316: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/$exit
      -- CP-element group 316: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_Update/ca
      -- CP-element group 316: 	 branch_block_stmt_436/assign_stmt_1547_to_assign_stmt_1557/type_cast_1550_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/$entry
      -- CP-element group 316: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/$entry
      -- CP-element group 316: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/$entry
      -- CP-element group 316: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/$entry
      -- CP-element group 316: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/$entry
      -- 
    ca_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1550_inst_ack_1, ack => convolution3D_CP_1120_elements(316)); -- 
    -- CP-element group 317:  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	426 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_Update/cr
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_Sample/ra
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_update_start_
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_sample_completed_
      -- 
    ra_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1588_inst_ack_0, ack => convolution3D_CP_1120_elements(317)); -- 
    cr_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(317), ack => RPIPE_maxpool_input_pipe_1588_inst_req_1); -- 
    -- CP-element group 318:  fork  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318: 	321 
    -- CP-element group 318:  members (9) 
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_Sample/rr
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_Sample/req
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_Update/ca
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_update_completed_
      -- 
    ca_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1588_inst_ack_1, ack => convolution3D_CP_1120_elements(318)); -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(318), ack => WPIPE_maxpool_output_pipe_1590_inst_req_0); -- 
    rr_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(318), ack => type_cast_1595_inst_req_0); -- 
    -- CP-element group 319:  transition  input  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (6) 
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_Update/req
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_Sample/ack
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_update_start_
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_sample_completed_
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1590_inst_ack_0, ack => convolution3D_CP_1120_elements(319)); -- 
    req_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(319), ack => WPIPE_maxpool_output_pipe_1590_inst_req_1); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	325 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_Update/ack
      -- CP-element group 320: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/WPIPE_maxpool_output_pipe_1590_update_completed_
      -- 
    ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1590_inst_ack_1, ack => convolution3D_CP_1120_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	318 
    -- CP-element group 321: successors 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_Sample/ra
      -- CP-element group 321: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_sample_completed_
      -- 
    ra_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1595_inst_ack_0, ack => convolution3D_CP_1120_elements(321)); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	426 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	325 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_Update/ca
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_update_completed_
      -- 
    ca_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1595_inst_ack_1, ack => convolution3D_CP_1120_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	426 
    -- CP-element group 323: successors 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_Sample/ra
      -- 
    ra_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1610_inst_ack_0, ack => convolution3D_CP_1120_elements(323)); -- 
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	426 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_Update/ca
      -- 
    ca_3427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1610_inst_ack_1, ack => convolution3D_CP_1120_elements(324)); -- 
    -- CP-element group 325:  branch  join  transition  place  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	320 
    -- CP-element group 325: 	322 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (10) 
      -- CP-element group 325: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616__exit__
      -- CP-element group 325: 	 branch_block_stmt_436/if_stmt_1617__entry__
      -- CP-element group 325: 	 branch_block_stmt_436/if_stmt_1617_dead_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_436/if_stmt_1617_eval_test/$entry
      -- CP-element group 325: 	 branch_block_stmt_436/if_stmt_1617_eval_test/$exit
      -- CP-element group 325: 	 branch_block_stmt_436/if_stmt_1617_eval_test/branch_req
      -- CP-element group 325: 	 branch_block_stmt_436/if_stmt_1617_if_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_436/if_stmt_1617_else_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_436/R_cmpx_xi428_1618_place
      -- CP-element group 325: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/$exit
      -- 
    branch_req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(325), ack => if_stmt_1617_branch_req_0); -- 
    convolution3D_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(320) & convolution3D_CP_1120_elements(322) & convolution3D_CP_1120_elements(324);
      gj_convolution3D_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  fork  transition  place  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	416 
    -- CP-element group 326: 	417 
    -- CP-element group 326: 	419 
    -- CP-element group 326: 	420 
    -- CP-element group 326:  members (20) 
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429
      -- CP-element group 326: 	 branch_block_stmt_436/if_stmt_1617_if_link/$exit
      -- CP-element group 326: 	 branch_block_stmt_436/if_stmt_1617_if_link/if_choice_transition
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/Update/cr
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1617_branch_ack_1, ack => convolution3D_CP_1120_elements(326)); -- 
    rr_4187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => type_cast_1566_inst_req_0); -- 
    cr_4192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => type_cast_1566_inst_req_1); -- 
    rr_4210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => type_cast_1573_inst_req_0); -- 
    cr_4215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => type_cast_1573_inst_req_1); -- 
    -- CP-element group 327:  fork  transition  place  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	427 
    -- CP-element group 327: 	428 
    -- CP-element group 327:  members (12) 
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437
      -- CP-element group 327: 	 branch_block_stmt_436/if_stmt_1617_else_link/else_choice_transition
      -- CP-element group 327: 	 branch_block_stmt_436/if_stmt_1617_else_link/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/rr
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1617_branch_ack_0, ack => convolution3D_CP_1120_elements(327)); -- 
    rr_4246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(327), ack => type_cast_1627_inst_req_0); -- 
    cr_4251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(327), ack => type_cast_1627_inst_req_1); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	430 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	334 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_Sample/ack
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_sample_complete
      -- 
    ack_3475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1656_index_offset_ack_0, ack => convolution3D_CP_1120_elements(328)); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	430 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (11) 
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_sample_start_
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_request/req
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_request/$entry
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_base_plus_offset/sum_rename_ack
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_base_plus_offset/sum_rename_req
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_base_plus_offset/$exit
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_base_plus_offset/$entry
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_Update/ack
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_offset_calculated
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_root_address_calculated
      -- 
    ack_3480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1656_index_offset_ack_1, ack => convolution3D_CP_1120_elements(329)); -- 
    req_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(329), ack => addr_of_1657_final_reg_req_0); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_request/ack
      -- CP-element group 330: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_request/$exit
      -- CP-element group 330: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_sample_completed_
      -- 
    ack_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1657_final_reg_ack_0, ack => convolution3D_CP_1120_elements(330)); -- 
    -- CP-element group 331:  join  fork  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	430 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (28) 
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_addr_resize/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_addr_resize/base_resize_req
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_addr_resize/base_resize_ack
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_plus_offset/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_plus_offset/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_plus_offset/sum_rename_req
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_addr_resize/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_address_resized
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_root_address_calculated
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_word_address_calculated
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_address_calculated
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_sample_start_
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_complete/ack
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/word_access_start/word_0/rr
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_complete/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/word_access_start/word_0/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/word_access_start/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/ptr_deref_1660_Split/split_ack
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/ptr_deref_1660_Split/split_req
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/ptr_deref_1660_Split/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/ptr_deref_1660_Split/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_word_addrgen/root_register_ack
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_word_addrgen/root_register_req
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_word_addrgen/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_word_addrgen/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_base_plus_offset/sum_rename_ack
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_update_completed_
      -- 
    ack_3495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1657_final_reg_ack_1, ack => convolution3D_CP_1120_elements(331)); -- 
    rr_3533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => ptr_deref_1660_store_0_req_0); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (5) 
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_sample_completed_
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/word_access_start/word_0/ra
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/word_access_start/word_0/$exit
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/word_access_start/$exit
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Sample/$exit
      -- 
    ra_3534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1660_store_0_ack_0, ack => convolution3D_CP_1120_elements(332)); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	430 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (5) 
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Update/word_access_complete/word_0/ca
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Update/word_access_complete/word_0/$exit
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_update_completed_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Update/word_access_complete/$exit
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Update/$exit
      -- 
    ca_3545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1660_store_0_ack_1, ack => convolution3D_CP_1120_elements(333)); -- 
    -- CP-element group 334:  join  transition  place  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	328 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	431 
    -- CP-element group 334:  members (5) 
      -- CP-element group 334: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662__exit__
      -- CP-element group 334: 	 branch_block_stmt_436/getRemainingElementsx_xexit437_ifx_xend353
      -- CP-element group 334: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/$exit
      -- CP-element group 334: 	 branch_block_stmt_436/getRemainingElementsx_xexit437_ifx_xend353_PhiReq/$entry
      -- CP-element group 334: 	 branch_block_stmt_436/getRemainingElementsx_xexit437_ifx_xend353_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(328) & convolution3D_CP_1120_elements(333);
      gj_convolution3D_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	431 
    -- CP-element group 335: successors 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_Sample/cra
      -- 
    cra_3557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1667_call_ack_0, ack => convolution3D_CP_1120_elements(335)); -- 
    -- CP-element group 336:  fork  transition  place  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	431 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336: 	339 
    -- CP-element group 336: 	343 
    -- CP-element group 336: 	344 
    -- CP-element group 336: 	345 
    -- CP-element group 336: 	346 
    -- CP-element group 336: 	347 
    -- CP-element group 336: 	348 
    -- CP-element group 336:  members (31) 
      -- CP-element group 336: 	 branch_block_stmt_436/call_stmt_1667__exit__
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735__entry__
      -- CP-element group 336: 	 branch_block_stmt_436/call_stmt_1667/$exit
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_Sample/rr
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_update_start_
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_Update/cr
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_Sample/rr
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_update_start_
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_Update/cr
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_Sample/rr
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_Sample/req
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_update_start_
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/$entry
      -- CP-element group 336: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_Update/cca
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_Update/cr
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_Sample/req
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_Update/$entry
      -- 
    cca_3562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1667_call_ack_1, ack => convolution3D_CP_1120_elements(336)); -- 
    rr_3615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(336), ack => type_cast_1710_inst_req_0); -- 
    cr_3648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(336), ack => type_cast_1729_inst_req_1); -- 
    rr_3643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(336), ack => type_cast_1729_inst_req_0); -- 
    cr_3634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(336), ack => type_cast_1720_inst_req_1); -- 
    rr_3629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(336), ack => type_cast_1720_inst_req_0); -- 
    req_3573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(336), ack => WPIPE_num_out_pipe_1679_inst_req_0); -- 
    cr_3620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(336), ack => type_cast_1710_inst_req_1); -- 
    req_3587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(336), ack => WPIPE_maxpool_output_pipe_1682_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_Update/req
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_update_start_
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_sample_completed_
      -- 
    ack_3574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1679_inst_ack_0, ack => convolution3D_CP_1120_elements(337)); -- 
    req_3578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(337), ack => WPIPE_num_out_pipe_1679_inst_req_1); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	349 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_num_out_pipe_1679_update_completed_
      -- 
    ack_3579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1679_inst_ack_1, ack => convolution3D_CP_1120_elements(338)); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	336 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_update_start_
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_Update/req
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_Sample/$exit
      -- 
    ack_3588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1682_inst_ack_0, ack => convolution3D_CP_1120_elements(339)); -- 
    req_3592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(339), ack => WPIPE_maxpool_output_pipe_1682_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_Sample/req
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1682_Update/$exit
      -- 
    ack_3593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1682_inst_ack_1, ack => convolution3D_CP_1120_elements(340)); -- 
    req_3601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(340), ack => WPIPE_maxpool_output_pipe_1686_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_Update/req
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_update_start_
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_sample_completed_
      -- 
    ack_3602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1686_inst_ack_0, ack => convolution3D_CP_1120_elements(341)); -- 
    req_3606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(341), ack => WPIPE_maxpool_output_pipe_1686_inst_req_1); -- 
    -- CP-element group 342:  transition  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	349 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/WPIPE_maxpool_output_pipe_1686_update_completed_
      -- 
    ack_3607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1686_inst_ack_1, ack => convolution3D_CP_1120_elements(342)); -- 
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	336 
    -- CP-element group 343: successors 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_Sample/ra
      -- CP-element group 343: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_sample_completed_
      -- 
    ra_3616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_0, ack => convolution3D_CP_1120_elements(343)); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	336 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	349 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_Update/ca
      -- CP-element group 344: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1710_Update/$exit
      -- 
    ca_3621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_1, ack => convolution3D_CP_1120_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	336 
    -- CP-element group 345: successors 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_Sample/ra
      -- CP-element group 345: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_sample_completed_
      -- 
    ra_3630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1720_inst_ack_0, ack => convolution3D_CP_1120_elements(345)); -- 
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	336 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	349 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_Update/ca
      -- CP-element group 346: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1720_update_completed_
      -- 
    ca_3635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1720_inst_ack_1, ack => convolution3D_CP_1120_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	336 
    -- CP-element group 347: successors 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_Sample/ra
      -- CP-element group 347: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_Sample/$exit
      -- 
    ra_3644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1729_inst_ack_0, ack => convolution3D_CP_1120_elements(347)); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	336 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_Update/ca
      -- CP-element group 348: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/type_cast_1729_update_completed_
      -- 
    ca_3649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1729_inst_ack_1, ack => convolution3D_CP_1120_elements(348)); -- 
    -- CP-element group 349:  join  transition  place  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	338 
    -- CP-element group 349: 	342 
    -- CP-element group 349: 	344 
    -- CP-element group 349: 	346 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	432 
    -- CP-element group 349:  members (6) 
      -- CP-element group 349: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735__exit__
      -- CP-element group 349: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody
      -- CP-element group 349: 	 branch_block_stmt_436/assign_stmt_1673_to_assign_stmt_1735/$exit
      -- CP-element group 349: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/$entry
      -- CP-element group 349: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1738/$entry
      -- CP-element group 349: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/$entry
      -- 
    convolution3D_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(338) & convolution3D_CP_1120_elements(342) & convolution3D_CP_1120_elements(344) & convolution3D_CP_1120_elements(346) & convolution3D_CP_1120_elements(348);
      gj_convolution3D_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	437 
    -- CP-element group 350: successors 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_sample_completed_
      -- CP-element group 350: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_Sample/ra
      -- CP-element group 350: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_Sample/$exit
      -- 
    ra_3661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1758_inst_ack_0, ack => convolution3D_CP_1120_elements(350)); -- 
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	437 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	354 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_Update/ca
      -- CP-element group 351: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_update_completed_
      -- CP-element group 351: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_Update/$exit
      -- 
    ca_3666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1758_inst_ack_1, ack => convolution3D_CP_1120_elements(351)); -- 
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	437 
    -- CP-element group 352: successors 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_Sample/ra
      -- 
    ra_3675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1762_inst_ack_0, ack => convolution3D_CP_1120_elements(352)); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	437 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_Update/ca
      -- 
    ca_3680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1762_inst_ack_1, ack => convolution3D_CP_1120_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	351 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_Sample/crr
      -- 
    crr_3688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(354), ack => call_stmt_1766_call_req_0); -- 
    convolution3D_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(351) & convolution3D_CP_1120_elements(353);
      gj_convolution3D_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_Sample/cra
      -- 
    cra_3689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1766_call_ack_0, ack => convolution3D_CP_1120_elements(355)); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	437 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	359 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_Update/cca
      -- 
    cca_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1766_call_ack_1, ack => convolution3D_CP_1120_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	437 
    -- CP-element group 357: successors 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_Sample/cra
      -- 
    cra_3703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1773_call_ack_0, ack => convolution3D_CP_1120_elements(357)); -- 
    -- CP-element group 358:  transition  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	437 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_Update/cca
      -- 
    cca_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1773_call_ack_1, ack => convolution3D_CP_1120_elements(358)); -- 
    -- CP-element group 359:  branch  join  transition  place  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	356 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (10) 
      -- CP-element group 359: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784__exit__
      -- CP-element group 359: 	 branch_block_stmt_436/if_stmt_1785__entry__
      -- CP-element group 359: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/$exit
      -- CP-element group 359: 	 branch_block_stmt_436/if_stmt_1785_dead_link/$entry
      -- CP-element group 359: 	 branch_block_stmt_436/if_stmt_1785_eval_test/$entry
      -- CP-element group 359: 	 branch_block_stmt_436/if_stmt_1785_eval_test/$exit
      -- CP-element group 359: 	 branch_block_stmt_436/if_stmt_1785_eval_test/branch_req
      -- CP-element group 359: 	 branch_block_stmt_436/R_exitcond5_1786_place
      -- CP-element group 359: 	 branch_block_stmt_436/if_stmt_1785_if_link/$entry
      -- CP-element group 359: 	 branch_block_stmt_436/if_stmt_1785_else_link/$entry
      -- 
    branch_req_3716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(359), ack => if_stmt_1785_branch_req_0); -- 
    convolution3D_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(356) & convolution3D_CP_1120_elements(358);
      gj_convolution3D_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	362 
    -- CP-element group 360: 	363 
    -- CP-element group 360:  members (18) 
      -- CP-element group 360: 	 branch_block_stmt_436/merge_stmt_1791__exit__
      -- CP-element group 360: 	 branch_block_stmt_436/assign_stmt_1796__entry__
      -- CP-element group 360: 	 branch_block_stmt_436/if_stmt_1785_if_link/$exit
      -- CP-element group 360: 	 branch_block_stmt_436/if_stmt_1785_if_link/if_choice_transition
      -- CP-element group 360: 	 branch_block_stmt_436/whilex_xbody_whilex_xend
      -- CP-element group 360: 	 branch_block_stmt_436/assign_stmt_1796/$entry
      -- CP-element group 360: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_update_start_
      -- CP-element group 360: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_Sample/rr
      -- CP-element group 360: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_Update/$entry
      -- CP-element group 360: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_Update/cr
      -- CP-element group 360: 	 branch_block_stmt_436/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 360: 	 branch_block_stmt_436/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 360: 	 branch_block_stmt_436/merge_stmt_1791_PhiReqMerge
      -- CP-element group 360: 	 branch_block_stmt_436/merge_stmt_1791_PhiAck/$entry
      -- CP-element group 360: 	 branch_block_stmt_436/merge_stmt_1791_PhiAck/$exit
      -- CP-element group 360: 	 branch_block_stmt_436/merge_stmt_1791_PhiAck/dummy
      -- 
    if_choice_transition_3721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1785_branch_ack_1, ack => convolution3D_CP_1120_elements(360)); -- 
    rr_3738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(360), ack => type_cast_1795_inst_req_0); -- 
    cr_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(360), ack => type_cast_1795_inst_req_1); -- 
    -- CP-element group 361:  fork  transition  place  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	433 
    -- CP-element group 361: 	434 
    -- CP-element group 361:  members (12) 
      -- CP-element group 361: 	 branch_block_stmt_436/if_stmt_1785_else_link/$exit
      -- CP-element group 361: 	 branch_block_stmt_436/if_stmt_1785_else_link/else_choice_transition
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/$entry
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/$entry
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/$entry
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/$entry
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/Sample/rr
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1785_branch_ack_0, ack => convolution3D_CP_1120_elements(361)); -- 
    rr_4299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(361), ack => type_cast_1741_inst_req_0); -- 
    cr_4304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(361), ack => type_cast_1741_inst_req_1); -- 
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: successors 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_sample_completed_
      -- CP-element group 362: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_Sample/ra
      -- 
    ra_3739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1795_inst_ack_0, ack => convolution3D_CP_1120_elements(362)); -- 
    -- CP-element group 363:  fork  transition  place  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	360 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363: 	365 
    -- CP-element group 363: 	367 
    -- CP-element group 363:  members (16) 
      -- CP-element group 363: 	 branch_block_stmt_436/assign_stmt_1796__exit__
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812__entry__
      -- CP-element group 363: 	 branch_block_stmt_436/assign_stmt_1796/$exit
      -- CP-element group 363: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_update_completed_
      -- CP-element group 363: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_436/assign_stmt_1796/type_cast_1795_Update/ca
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/$entry
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_update_start_
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_Sample/crr
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_Update/ccr
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_update_start_
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_Update/cr
      -- 
    ca_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1795_inst_ack_1, ack => convolution3D_CP_1120_elements(363)); -- 
    crr_3755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(363), ack => call_stmt_1799_call_req_0); -- 
    ccr_3760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(363), ack => call_stmt_1799_call_req_1); -- 
    cr_3774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(363), ack => type_cast_1803_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_sample_completed_
      -- CP-element group 364: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_Sample/cra
      -- 
    cra_3756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1799_call_ack_0, ack => convolution3D_CP_1120_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_update_completed_
      -- CP-element group 365: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/call_stmt_1799_Update/cca
      -- CP-element group 365: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_Sample/rr
      -- 
    cca_3761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1799_call_ack_1, ack => convolution3D_CP_1120_elements(365)); -- 
    rr_3769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(365), ack => type_cast_1803_inst_req_0); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_Sample/ra
      -- 
    ra_3770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1803_inst_ack_0, ack => convolution3D_CP_1120_elements(366)); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	363 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/type_cast_1803_Update/ca
      -- CP-element group 367: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_sample_start_
      -- CP-element group 367: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_Sample/req
      -- 
    ca_3775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1803_inst_ack_1, ack => convolution3D_CP_1120_elements(367)); -- 
    req_3783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(367), ack => WPIPE_elapsed_time_pipe_1810_inst_req_0); -- 
    -- CP-element group 368:  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_Sample/ack
      -- CP-element group 368: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_Update/req
      -- 
    ack_3784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1810_inst_ack_0, ack => convolution3D_CP_1120_elements(368)); -- 
    req_3788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => WPIPE_elapsed_time_pipe_1810_inst_req_1); -- 
    -- CP-element group 369:  transition  place  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369:  members (16) 
      -- CP-element group 369: 	 $exit
      -- CP-element group 369: 	 branch_block_stmt_436/$exit
      -- CP-element group 369: 	 branch_block_stmt_436/branch_block_stmt_436__exit__
      -- CP-element group 369: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812__exit__
      -- CP-element group 369: 	 branch_block_stmt_436/return__
      -- CP-element group 369: 	 branch_block_stmt_436/merge_stmt_1815__exit__
      -- CP-element group 369: 	 branch_block_stmt_436/merge_stmt_1815_PhiReqMerge
      -- CP-element group 369: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/$exit
      -- CP-element group 369: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_436/call_stmt_1799_to_assign_stmt_1812/WPIPE_elapsed_time_pipe_1810_Update/ack
      -- CP-element group 369: 	 branch_block_stmt_436/return___PhiReq/$entry
      -- CP-element group 369: 	 branch_block_stmt_436/return___PhiReq/$exit
      -- CP-element group 369: 	 branch_block_stmt_436/merge_stmt_1815_PhiAck/$entry
      -- CP-element group 369: 	 branch_block_stmt_436/merge_stmt_1815_PhiAck/$exit
      -- CP-element group 369: 	 branch_block_stmt_436/merge_stmt_1815_PhiAck/dummy
      -- 
    ack_3789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1810_inst_ack_1, ack => convolution3D_CP_1120_elements(369)); -- 
    -- CP-element group 370:  transition  output  delay-element  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	138 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	374 
    -- CP-element group 370:  members (5) 
      -- CP-element group 370: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/$exit
      -- CP-element group 370: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_801/$exit
      -- CP-element group 370: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/$exit
      -- CP-element group 370: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_805_konst_delay_trans
      -- CP-element group 370: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_req
      -- 
    phi_stmt_801_req_3812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_801_req_3812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(370), ack => phi_stmt_801_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(370) is a control-delay.
    cp_element_370_delay: control_delay_element  generic map(name => " 370_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(138), ack => convolution3D_CP_1120_elements(370), clk => clk, reset =>reset);
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	203 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	373 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/Sample/ra
      -- 
    ra_3832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_0, ack => convolution3D_CP_1120_elements(371)); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	203 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (2) 
      -- CP-element group 372: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/Update/ca
      -- 
    ca_3837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_1, ack => convolution3D_CP_1120_elements(372)); -- 
    -- CP-element group 373:  join  transition  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	371 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (6) 
      -- CP-element group 373: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 373: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/$exit
      -- CP-element group 373: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/$exit
      -- CP-element group 373: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/$exit
      -- CP-element group 373: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_sources/type_cast_807/SplitProtocol/$exit
      -- CP-element group 373: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_801/phi_stmt_801_req
      -- 
    phi_stmt_801_req_3838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_801_req_3838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(373), ack => phi_stmt_801_req_1); -- 
    convolution3D_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(371) & convolution3D_CP_1120_elements(372);
      gj_convolution3D_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  merge  transition  place  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: 	370 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (2) 
      -- CP-element group 374: 	 branch_block_stmt_436/merge_stmt_800_PhiReqMerge
      -- CP-element group 374: 	 branch_block_stmt_436/merge_stmt_800_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(374) <= OrReduce(convolution3D_CP_1120_elements(373) & convolution3D_CP_1120_elements(370));
    -- CP-element group 375:  fork  transition  place  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	139 
    -- CP-element group 375: 	140 
    -- CP-element group 375: 	142 
    -- CP-element group 375: 	143 
    -- CP-element group 375: 	148 
    -- CP-element group 375: 	155 
    -- CP-element group 375: 	162 
    -- CP-element group 375: 	169 
    -- CP-element group 375: 	176 
    -- CP-element group 375: 	183 
    -- CP-element group 375: 	190 
    -- CP-element group 375: 	197 
    -- CP-element group 375: 	200 
    -- CP-element group 375:  members (56) 
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Update/word_access_complete/word_0/cr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Update/word_access_complete/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Update/word_access_complete/word_0/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/merge_stmt_800__exit__
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987__entry__
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_Update/cr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/ptr_deref_974_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_945_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_Update/cr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_966_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_resized_1
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_scaled_1
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_computed_1
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_resize_1/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_resize_1/$exit
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_resize_1/index_resize_req
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_resize_1/index_resize_ack
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_scale_1/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_scale_1/$exit
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_scale_1/scale_rename_req
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_index_scale_1/scale_rename_ack
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_update_start
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_Sample/req
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/array_obj_ref_813_final_index_sum_regn_Update/req
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_complete/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/addr_of_814_complete/req
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/RPIPE_maxpool_input_pipe_817_Sample/rr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_824_Update/cr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_840_Update/cr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_861_Update/cr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_882_Update/cr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_903_Update/cr
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_update_start_
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_436/assign_stmt_815_to_assign_stmt_987/type_cast_924_Update/cr
      -- CP-element group 375: 	 branch_block_stmt_436/merge_stmt_800_PhiAck/$exit
      -- CP-element group 375: 	 branch_block_stmt_436/merge_stmt_800_PhiAck/phi_stmt_801_ack
      -- 
    phi_stmt_801_ack_3843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_801_ack_0, ack => convolution3D_CP_1120_elements(375)); -- 
    cr_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => ptr_deref_974_store_0_req_1); -- 
    cr_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => type_cast_945_inst_req_1); -- 
    cr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => type_cast_966_inst_req_1); -- 
    req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => array_obj_ref_813_index_offset_req_0); -- 
    req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => array_obj_ref_813_index_offset_req_1); -- 
    req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => addr_of_814_final_reg_req_1); -- 
    rr_2105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => RPIPE_maxpool_input_pipe_817_inst_req_0); -- 
    cr_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => type_cast_824_inst_req_1); -- 
    cr_2180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => type_cast_840_inst_req_1); -- 
    cr_2222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => type_cast_861_inst_req_1); -- 
    cr_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => type_cast_882_inst_req_1); -- 
    cr_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => type_cast_903_inst_req_1); -- 
    cr_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => type_cast_924_inst_req_1); -- 
    -- CP-element group 376:  transition  output  delay-element  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	128 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	380 
    -- CP-element group 376:  members (5) 
      -- CP-element group 376: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/$exit
      -- CP-element group 376: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1019/$exit
      -- CP-element group 376: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/$exit
      -- CP-element group 376: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1025_konst_delay_trans
      -- CP-element group 376: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_req
      -- 
    phi_stmt_1019_req_3866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1019_req_3866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(376), ack => phi_stmt_1019_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(376) is a control-delay.
    cp_element_376_delay: control_delay_element  generic map(name => " 376_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(128), ack => convolution3D_CP_1120_elements(376), clk => clk, reset =>reset);
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	202 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (2) 
      -- CP-element group 377: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/Sample/ra
      -- 
    ra_3886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1022_inst_ack_0, ack => convolution3D_CP_1120_elements(377)); -- 
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	202 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (2) 
      -- CP-element group 378: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/Update/ca
      -- 
    ca_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1022_inst_ack_1, ack => convolution3D_CP_1120_elements(378)); -- 
    -- CP-element group 379:  join  transition  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (6) 
      -- CP-element group 379: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 379: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/$exit
      -- CP-element group 379: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/$exit
      -- CP-element group 379: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/$exit
      -- CP-element group 379: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_sources/type_cast_1022/SplitProtocol/$exit
      -- CP-element group 379: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1019/phi_stmt_1019_req
      -- 
    phi_stmt_1019_req_3892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1019_req_3892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(379), ack => phi_stmt_1019_req_0); -- 
    convolution3D_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(377) & convolution3D_CP_1120_elements(378);
      gj_convolution3D_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  merge  transition  place  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	376 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (2) 
      -- CP-element group 380: 	 branch_block_stmt_436/merge_stmt_1018_PhiReqMerge
      -- CP-element group 380: 	 branch_block_stmt_436/merge_stmt_1018_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(380) <= OrReduce(convolution3D_CP_1120_elements(376) & convolution3D_CP_1120_elements(379));
    -- CP-element group 381:  branch  transition  place  input  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	204 
    -- CP-element group 381: 	205 
    -- CP-element group 381:  members (15) 
      -- CP-element group 381: 	 branch_block_stmt_436/merge_stmt_1018__exit__
      -- CP-element group 381: 	 branch_block_stmt_436/assign_stmt_1032_to_assign_stmt_1038__entry__
      -- CP-element group 381: 	 branch_block_stmt_436/assign_stmt_1032_to_assign_stmt_1038__exit__
      -- CP-element group 381: 	 branch_block_stmt_436/if_stmt_1039__entry__
      -- CP-element group 381: 	 branch_block_stmt_436/if_stmt_1039_else_link/$entry
      -- CP-element group 381: 	 branch_block_stmt_436/if_stmt_1039_if_link/$entry
      -- CP-element group 381: 	 branch_block_stmt_436/if_stmt_1039_eval_test/branch_req
      -- CP-element group 381: 	 branch_block_stmt_436/if_stmt_1039_eval_test/$exit
      -- CP-element group 381: 	 branch_block_stmt_436/if_stmt_1039_eval_test/$entry
      -- CP-element group 381: 	 branch_block_stmt_436/if_stmt_1039_dead_link/$entry
      -- CP-element group 381: 	 branch_block_stmt_436/assign_stmt_1032_to_assign_stmt_1038/$exit
      -- CP-element group 381: 	 branch_block_stmt_436/assign_stmt_1032_to_assign_stmt_1038/$entry
      -- CP-element group 381: 	 branch_block_stmt_436/R_tobool_1040_place
      -- CP-element group 381: 	 branch_block_stmt_436/merge_stmt_1018_PhiAck/$exit
      -- CP-element group 381: 	 branch_block_stmt_436/merge_stmt_1018_PhiAck/phi_stmt_1019_ack
      -- 
    phi_stmt_1019_ack_3897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1019_ack_0, ack => convolution3D_CP_1120_elements(381)); -- 
    branch_req_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(381), ack => if_stmt_1039_branch_req_0); -- 
    -- CP-element group 382:  transition  output  delay-element  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	205 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	384 
    -- CP-element group 382:  members (4) 
      -- CP-element group 382: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/$exit
      -- CP-element group 382: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/$exit
      -- CP-element group 382: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1064_konst_delay_trans
      -- CP-element group 382: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_req
      -- 
    phi_stmt_1060_req_3920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1060_req_3920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(382), ack => phi_stmt_1060_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(382) is a control-delay.
    cp_element_382_delay: control_delay_element  generic map(name => " 382_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(205), ack => convolution3D_CP_1120_elements(382), clk => clk, reset =>reset);
    -- CP-element group 383:  transition  output  delay-element  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	205 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (4) 
      -- CP-element group 383: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/$exit
      -- CP-element group 383: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/$exit
      -- CP-element group 383: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1071_konst_delay_trans
      -- CP-element group 383: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_req
      -- 
    phi_stmt_1067_req_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1067_req_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(383), ack => phi_stmt_1067_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(383) is a control-delay.
    cp_element_383_delay: control_delay_element  generic map(name => " 383_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(205), ack => convolution3D_CP_1120_elements(383), clk => clk, reset =>reset);
    -- CP-element group 384:  join  transition  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	382 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	392 
    -- CP-element group 384:  members (1) 
      -- CP-element group 384: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(382) & convolution3D_CP_1120_elements(383);
      gj_convolution3D_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	215 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (2) 
      -- CP-element group 385: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/Sample/ra
      -- 
    ra_3948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1066_inst_ack_0, ack => convolution3D_CP_1120_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	215 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (2) 
      -- CP-element group 386: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/Update/ca
      -- 
    ca_3953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1066_inst_ack_1, ack => convolution3D_CP_1120_elements(386)); -- 
    -- CP-element group 387:  join  transition  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	391 
    -- CP-element group 387:  members (5) 
      -- CP-element group 387: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/$exit
      -- CP-element group 387: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/$exit
      -- CP-element group 387: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/$exit
      -- CP-element group 387: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1066/SplitProtocol/$exit
      -- CP-element group 387: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1060/phi_stmt_1060_req
      -- 
    phi_stmt_1060_req_3954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1060_req_3954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(387), ack => phi_stmt_1060_req_1); -- 
    convolution3D_cp_element_group_387: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_387"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(385) & convolution3D_CP_1120_elements(386);
      gj_convolution3D_cp_element_group_387 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(387), clk => clk, reset => reset); --
    end block;
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	215 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	390 
    -- CP-element group 388:  members (2) 
      -- CP-element group 388: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/Sample/ra
      -- 
    ra_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_0, ack => convolution3D_CP_1120_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	215 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (2) 
      -- CP-element group 389: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/Update/ca
      -- 
    ca_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_1, ack => convolution3D_CP_1120_elements(389)); -- 
    -- CP-element group 390:  join  transition  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	388 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (5) 
      -- CP-element group 390: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/$exit
      -- CP-element group 390: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/$exit
      -- CP-element group 390: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/$exit
      -- CP-element group 390: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_sources/type_cast_1073/SplitProtocol/$exit
      -- CP-element group 390: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1067/phi_stmt_1067_req
      -- 
    phi_stmt_1067_req_3977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1067_req_3977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(390), ack => phi_stmt_1067_req_1); -- 
    convolution3D_cp_element_group_390: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_390"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(388) & convolution3D_CP_1120_elements(389);
      gj_convolution3D_cp_element_group_390 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(390), clk => clk, reset => reset); --
    end block;
    -- CP-element group 391:  join  transition  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	387 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (1) 
      -- CP-element group 391: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(387) & convolution3D_CP_1120_elements(390);
      gj_convolution3D_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  merge  fork  transition  place  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: 	384 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392: 	394 
    -- CP-element group 392:  members (2) 
      -- CP-element group 392: 	 branch_block_stmt_436/merge_stmt_1059_PhiReqMerge
      -- CP-element group 392: 	 branch_block_stmt_436/merge_stmt_1059_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(392) <= OrReduce(convolution3D_CP_1120_elements(391) & convolution3D_CP_1120_elements(384));
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	395 
    -- CP-element group 393:  members (1) 
      -- CP-element group 393: 	 branch_block_stmt_436/merge_stmt_1059_PhiAck/phi_stmt_1060_ack
      -- 
    phi_stmt_1060_ack_3982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1060_ack_0, ack => convolution3D_CP_1120_elements(393)); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	392 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (1) 
      -- CP-element group 394: 	 branch_block_stmt_436/merge_stmt_1059_PhiAck/phi_stmt_1067_ack
      -- 
    phi_stmt_1067_ack_3983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1067_ack_0, ack => convolution3D_CP_1120_elements(394)); -- 
    -- CP-element group 395:  join  fork  transition  place  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	393 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	206 
    -- CP-element group 395: 	211 
    -- CP-element group 395: 	212 
    -- CP-element group 395: 	213 
    -- CP-element group 395:  members (16) 
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_sample_start_
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_update_start_
      -- CP-element group 395: 	 branch_block_stmt_436/merge_stmt_1059__exit__
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116__entry__
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_Sample/$entry
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_Sample/rr
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_Sample/$entry
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_Update/cr
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/RPIPE_maxpool_input_pipe_1088_sample_start_
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/$entry
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_Update/cr
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1110_Sample/rr
      -- CP-element group 395: 	 branch_block_stmt_436/assign_stmt_1080_to_assign_stmt_1116/type_cast_1095_update_start_
      -- CP-element group 395: 	 branch_block_stmt_436/merge_stmt_1059_PhiAck/$exit
      -- 
    rr_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(395), ack => RPIPE_maxpool_input_pipe_1088_inst_req_0); -- 
    cr_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(395), ack => type_cast_1095_inst_req_1); -- 
    cr_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(395), ack => type_cast_1110_inst_req_1); -- 
    rr_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(395), ack => type_cast_1110_inst_req_0); -- 
    convolution3D_cp_element_group_395: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_395"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(393) & convolution3D_CP_1120_elements(394);
      gj_convolution3D_cp_element_group_395 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(395), clk => clk, reset => reset); --
    end block;
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	216 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	398 
    -- CP-element group 396:  members (2) 
      -- CP-element group 396: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/Sample/ra
      -- 
    ra_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1127_inst_ack_0, ack => convolution3D_CP_1120_elements(396)); -- 
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	216 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (2) 
      -- CP-element group 397: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/Update/ca
      -- 
    ca_4012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1127_inst_ack_1, ack => convolution3D_CP_1120_elements(397)); -- 
    -- CP-element group 398:  join  transition  place  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	396 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (8) 
      -- CP-element group 398: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 398: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/$exit
      -- CP-element group 398: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/$exit
      -- CP-element group 398: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/$exit
      -- CP-element group 398: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_sources/type_cast_1127/SplitProtocol/$exit
      -- CP-element group 398: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1124/phi_stmt_1124_req
      -- CP-element group 398: 	 branch_block_stmt_436/merge_stmt_1123_PhiReqMerge
      -- CP-element group 398: 	 branch_block_stmt_436/merge_stmt_1123_PhiAck/$entry
      -- 
    phi_stmt_1124_req_4013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1124_req_4013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(398), ack => phi_stmt_1124_req_0); -- 
    convolution3D_cp_element_group_398: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_398"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(396) & convolution3D_CP_1120_elements(397);
      gj_convolution3D_cp_element_group_398 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(398), clk => clk, reset => reset); --
    end block;
    -- CP-element group 399:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	217 
    -- CP-element group 399: 	218 
    -- CP-element group 399: 	220 
    -- CP-element group 399: 	222 
    -- CP-element group 399:  members (29) 
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_scale_1/scale_rename_ack
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_scale_1/scale_rename_req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Update/word_access_complete/word_0/cr
      -- CP-element group 399: 	 branch_block_stmt_436/merge_stmt_1123__exit__
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162__entry__
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_update_start
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_resized_1
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_scale_1/$exit
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Update/word_access_complete/word_0/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_scale_1/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Update/word_access_complete/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/ptr_deref_1160_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_complete/req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/addr_of_1157_complete/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_resize_1/index_resize_ack
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_resize_1/index_resize_req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_resize_1/$exit
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_resize_1/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_computed_1
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_index_scaled_1
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_Update/req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1134_to_assign_stmt_1162/array_obj_ref_1156_final_index_sum_regn_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/merge_stmt_1123_PhiAck/$exit
      -- CP-element group 399: 	 branch_block_stmt_436/merge_stmt_1123_PhiAck/phi_stmt_1124_ack
      -- 
    phi_stmt_1124_ack_4018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1124_ack_0, ack => convolution3D_CP_1120_elements(399)); -- 
    cr_2706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => ptr_deref_1160_store_0_req_1); -- 
    req_2656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => addr_of_1157_final_reg_req_1); -- 
    req_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => array_obj_ref_1156_index_offset_req_1); -- 
    req_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => array_obj_ref_1156_index_offset_req_0); -- 
    -- CP-element group 400:  merge  fork  transition  place  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	204 
    -- CP-element group 400: 	223 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	224 
    -- CP-element group 400: 	225 
    -- CP-element group 400: 	226 
    -- CP-element group 400: 	227 
    -- CP-element group 400: 	228 
    -- CP-element group 400: 	229 
    -- CP-element group 400: 	230 
    -- CP-element group 400: 	231 
    -- CP-element group 400:  members (31) 
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_update_start_
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_sample_start_
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_Update/cr
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_update_start_
      -- CP-element group 400: 	 branch_block_stmt_436/merge_stmt_1164__exit__
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216__entry__
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_sample_start_
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_Sample/rr
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1167_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_Sample/rr
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1171_Update/cr
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_sample_start_
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_update_start_
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_Sample/rr
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1175_Update/cr
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_sample_start_
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_update_start_
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_Sample/rr
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/assign_stmt_1168_to_assign_stmt_1216/type_cast_1179_Update/cr
      -- CP-element group 400: 	 branch_block_stmt_436/merge_stmt_1164_PhiReqMerge
      -- CP-element group 400: 	 branch_block_stmt_436/merge_stmt_1164_PhiAck/$entry
      -- CP-element group 400: 	 branch_block_stmt_436/merge_stmt_1164_PhiAck/$exit
      -- CP-element group 400: 	 branch_block_stmt_436/merge_stmt_1164_PhiAck/dummy
      -- 
    cr_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(400), ack => type_cast_1167_inst_req_1); -- 
    rr_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(400), ack => type_cast_1167_inst_req_0); -- 
    rr_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(400), ack => type_cast_1171_inst_req_0); -- 
    cr_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(400), ack => type_cast_1171_inst_req_1); -- 
    rr_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(400), ack => type_cast_1175_inst_req_0); -- 
    cr_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(400), ack => type_cast_1175_inst_req_1); -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(400), ack => type_cast_1179_inst_req_0); -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(400), ack => type_cast_1179_inst_req_1); -- 
    convolution3D_CP_1120_elements(400) <= OrReduce(convolution3D_CP_1120_elements(204) & convolution3D_CP_1120_elements(223));
    -- CP-element group 401:  transition  output  delay-element  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	247 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	405 
    -- CP-element group 401:  members (5) 
      -- CP-element group 401: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/$exit
      -- CP-element group 401: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1297/$exit
      -- CP-element group 401: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/$exit
      -- CP-element group 401: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1301_konst_delay_trans
      -- CP-element group 401: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_req
      -- 
    phi_stmt_1297_req_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1297_req_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(401), ack => phi_stmt_1297_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(401) is a control-delay.
    cp_element_401_delay: control_delay_element  generic map(name => " 401_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(247), ack => convolution3D_CP_1120_elements(401), clk => clk, reset =>reset);
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	312 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (2) 
      -- CP-element group 402: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Sample/$exit
      -- CP-element group 402: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Sample/ra
      -- 
    ra_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1303_inst_ack_0, ack => convolution3D_CP_1120_elements(402)); -- 
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	312 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (2) 
      -- CP-element group 403: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Update/$exit
      -- CP-element group 403: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Update/ca
      -- 
    ca_4077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1303_inst_ack_1, ack => convolution3D_CP_1120_elements(403)); -- 
    -- CP-element group 404:  join  transition  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (6) 
      -- CP-element group 404: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/$exit
      -- CP-element group 404: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/$exit
      -- CP-element group 404: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/$exit
      -- CP-element group 404: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/$exit
      -- CP-element group 404: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/$exit
      -- CP-element group 404: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1297/phi_stmt_1297_req
      -- 
    phi_stmt_1297_req_4078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1297_req_4078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(404), ack => phi_stmt_1297_req_1); -- 
    convolution3D_cp_element_group_404: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_404"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(402) & convolution3D_CP_1120_elements(403);
      gj_convolution3D_cp_element_group_404 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(404), clk => clk, reset => reset); --
    end block;
    -- CP-element group 405:  merge  transition  place  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	401 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (2) 
      -- CP-element group 405: 	 branch_block_stmt_436/merge_stmt_1296_PhiReqMerge
      -- CP-element group 405: 	 branch_block_stmt_436/merge_stmt_1296_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(405) <= OrReduce(convolution3D_CP_1120_elements(401) & convolution3D_CP_1120_elements(404));
    -- CP-element group 406:  fork  transition  place  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	292 
    -- CP-element group 406: 	309 
    -- CP-element group 406: 	306 
    -- CP-element group 406: 	299 
    -- CP-element group 406: 	248 
    -- CP-element group 406: 	249 
    -- CP-element group 406: 	251 
    -- CP-element group 406: 	252 
    -- CP-element group 406: 	257 
    -- CP-element group 406: 	264 
    -- CP-element group 406: 	271 
    -- CP-element group 406: 	278 
    -- CP-element group 406: 	285 
    -- CP-element group 406:  members (56) 
      -- CP-element group 406: 	 branch_block_stmt_436/merge_stmt_1296__exit__
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483__entry__
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_resized_1
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_scaled_1
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_computed_1
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Update/word_access_complete/word_0/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_resize_1/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_resize_1/$exit
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_resize_1/index_resize_req
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_resize_1/index_resize_ack
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_scale_1/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_scale_1/$exit
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_scale_1/scale_rename_req
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_index_scale_1/scale_rename_ack
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_update_start
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_Sample/req
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/array_obj_ref_1309_final_index_sum_regn_Update/req
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Update/word_access_complete/word_0/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_Update/word_access_complete/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_complete/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/addr_of_1310_complete/req
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/RPIPE_maxpool_input_pipe_1313_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1320_Update/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1336_Update/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1357_Update/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1378_Update/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1399_Update/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1420_Update/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1441_Update/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/type_cast_1462_Update/cr
      -- CP-element group 406: 	 branch_block_stmt_436/assign_stmt_1311_to_assign_stmt_1483/ptr_deref_1470_update_start_
      -- CP-element group 406: 	 branch_block_stmt_436/merge_stmt_1296_PhiAck/$exit
      -- CP-element group 406: 	 branch_block_stmt_436/merge_stmt_1296_PhiAck/phi_stmt_1297_ack
      -- 
    phi_stmt_1297_ack_4083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1297_ack_0, ack => convolution3D_CP_1120_elements(406)); -- 
    cr_3306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => ptr_deref_1470_store_0_req_1); -- 
    req_2900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => array_obj_ref_1309_index_offset_req_0); -- 
    req_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => array_obj_ref_1309_index_offset_req_1); -- 
    req_2920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => addr_of_1310_final_reg_req_1); -- 
    rr_2929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => RPIPE_maxpool_input_pipe_1313_inst_req_0); -- 
    cr_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => type_cast_1320_inst_req_1); -- 
    cr_3004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => type_cast_1336_inst_req_1); -- 
    cr_3046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => type_cast_1357_inst_req_1); -- 
    cr_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => type_cast_1378_inst_req_1); -- 
    cr_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => type_cast_1399_inst_req_1); -- 
    cr_3172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => type_cast_1420_inst_req_1); -- 
    cr_3214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => type_cast_1441_inst_req_1); -- 
    cr_3256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => type_cast_1462_inst_req_1); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	311 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	409 
    -- CP-element group 407:  members (2) 
      -- CP-element group 407: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/ra
      -- 
    ra_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_0, ack => convolution3D_CP_1120_elements(407)); -- 
    -- CP-element group 408:  transition  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	311 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (2) 
      -- CP-element group 408: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/ca
      -- 
    ca_4120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_1, ack => convolution3D_CP_1120_elements(408)); -- 
    -- CP-element group 409:  join  transition  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	407 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	411 
    -- CP-element group 409:  members (6) 
      -- CP-element group 409: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/$exit
      -- CP-element group 409: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/$exit
      -- CP-element group 409: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$exit
      -- CP-element group 409: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/$exit
      -- CP-element group 409: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/$exit
      -- CP-element group 409: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_req
      -- 
    phi_stmt_1515_req_4121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_req_4121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(409), ack => phi_stmt_1515_req_1); -- 
    convolution3D_cp_element_group_409: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_409"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(407) & convolution3D_CP_1120_elements(408);
      gj_convolution3D_cp_element_group_409 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(409), clk => clk, reset => reset); --
    end block;
    -- CP-element group 410:  transition  output  delay-element  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	234 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (5) 
      -- CP-element group 410: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/$exit
      -- CP-element group 410: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1515/$exit
      -- CP-element group 410: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$exit
      -- CP-element group 410: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1519_konst_delay_trans
      -- CP-element group 410: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1515/phi_stmt_1515_req
      -- 
    phi_stmt_1515_req_4132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_req_4132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(410), ack => phi_stmt_1515_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(410) is a control-delay.
    cp_element_410_delay: control_delay_element  generic map(name => " 410_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(234), ack => convolution3D_CP_1120_elements(410), clk => clk, reset =>reset);
    -- CP-element group 411:  merge  transition  place  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: 	409 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (2) 
      -- CP-element group 411: 	 branch_block_stmt_436/merge_stmt_1514_PhiReqMerge
      -- CP-element group 411: 	 branch_block_stmt_436/merge_stmt_1514_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(411) <= OrReduce(convolution3D_CP_1120_elements(410) & convolution3D_CP_1120_elements(409));
    -- CP-element group 412:  branch  transition  place  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	313 
    -- CP-element group 412: 	314 
    -- CP-element group 412:  members (15) 
      -- CP-element group 412: 	 branch_block_stmt_436/merge_stmt_1514__exit__
      -- CP-element group 412: 	 branch_block_stmt_436/assign_stmt_1528_to_assign_stmt_1534__entry__
      -- CP-element group 412: 	 branch_block_stmt_436/assign_stmt_1528_to_assign_stmt_1534__exit__
      -- CP-element group 412: 	 branch_block_stmt_436/if_stmt_1535__entry__
      -- CP-element group 412: 	 branch_block_stmt_436/R_tobool344_1536_place
      -- CP-element group 412: 	 branch_block_stmt_436/if_stmt_1535_else_link/$entry
      -- CP-element group 412: 	 branch_block_stmt_436/if_stmt_1535_if_link/$entry
      -- CP-element group 412: 	 branch_block_stmt_436/if_stmt_1535_eval_test/branch_req
      -- CP-element group 412: 	 branch_block_stmt_436/if_stmt_1535_eval_test/$exit
      -- CP-element group 412: 	 branch_block_stmt_436/if_stmt_1535_eval_test/$entry
      -- CP-element group 412: 	 branch_block_stmt_436/if_stmt_1535_dead_link/$entry
      -- CP-element group 412: 	 branch_block_stmt_436/assign_stmt_1528_to_assign_stmt_1534/$exit
      -- CP-element group 412: 	 branch_block_stmt_436/assign_stmt_1528_to_assign_stmt_1534/$entry
      -- CP-element group 412: 	 branch_block_stmt_436/merge_stmt_1514_PhiAck/$exit
      -- CP-element group 412: 	 branch_block_stmt_436/merge_stmt_1514_PhiAck/phi_stmt_1515_ack
      -- 
    phi_stmt_1515_ack_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1515_ack_0, ack => convolution3D_CP_1120_elements(412)); -- 
    branch_req_3340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(412), ack => if_stmt_1535_branch_req_0); -- 
    -- CP-element group 413:  transition  output  delay-element  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	316 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	415 
    -- CP-element group 413:  members (4) 
      -- CP-element group 413: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/$exit
      -- CP-element group 413: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/$exit
      -- CP-element group 413: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1564_konst_delay_trans
      -- CP-element group 413: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_req
      -- 
    phi_stmt_1560_req_4160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1560_req_4160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(413), ack => phi_stmt_1560_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(413) is a control-delay.
    cp_element_413_delay: control_delay_element  generic map(name => " 413_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(316), ack => convolution3D_CP_1120_elements(413), clk => clk, reset =>reset);
    -- CP-element group 414:  transition  output  delay-element  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	316 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (4) 
      -- CP-element group 414: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/$exit
      -- CP-element group 414: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/$exit
      -- CP-element group 414: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1571_konst_delay_trans
      -- CP-element group 414: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_req
      -- 
    phi_stmt_1567_req_4168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1567_req_4168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(414), ack => phi_stmt_1567_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(414) is a control-delay.
    cp_element_414_delay: control_delay_element  generic map(name => " 414_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(316), ack => convolution3D_CP_1120_elements(414), clk => clk, reset =>reset);
    -- CP-element group 415:  join  transition  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: 	413 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	423 
    -- CP-element group 415:  members (1) 
      -- CP-element group 415: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(414) & convolution3D_CP_1120_elements(413);
      gj_convolution3D_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  transition  input  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	326 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	418 
    -- CP-element group 416:  members (2) 
      -- CP-element group 416: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/Sample/ra
      -- 
    ra_4188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1566_inst_ack_0, ack => convolution3D_CP_1120_elements(416)); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	326 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (2) 
      -- CP-element group 417: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/Update/ca
      -- 
    ca_4193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1566_inst_ack_1, ack => convolution3D_CP_1120_elements(417)); -- 
    -- CP-element group 418:  join  transition  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	416 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	422 
    -- CP-element group 418:  members (5) 
      -- CP-element group 418: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/$exit
      -- CP-element group 418: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/$exit
      -- CP-element group 418: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/$exit
      -- CP-element group 418: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_sources/type_cast_1566/SplitProtocol/$exit
      -- CP-element group 418: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1560/phi_stmt_1560_req
      -- 
    phi_stmt_1560_req_4194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1560_req_4194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(418), ack => phi_stmt_1560_req_1); -- 
    convolution3D_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(416) & convolution3D_CP_1120_elements(417);
      gj_convolution3D_cp_element_group_418 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	326 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	421 
    -- CP-element group 419:  members (2) 
      -- CP-element group 419: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/Sample/ra
      -- 
    ra_4211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1573_inst_ack_0, ack => convolution3D_CP_1120_elements(419)); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	326 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (2) 
      -- CP-element group 420: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/Update/ca
      -- 
    ca_4216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1573_inst_ack_1, ack => convolution3D_CP_1120_elements(420)); -- 
    -- CP-element group 421:  join  transition  output  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	419 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (5) 
      -- CP-element group 421: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/$exit
      -- CP-element group 421: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/$exit
      -- CP-element group 421: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/$exit
      -- CP-element group 421: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_sources/type_cast_1573/SplitProtocol/$exit
      -- CP-element group 421: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1567/phi_stmt_1567_req
      -- 
    phi_stmt_1567_req_4217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1567_req_4217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(421), ack => phi_stmt_1567_req_1); -- 
    convolution3D_cp_element_group_421: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_421"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(419) & convolution3D_CP_1120_elements(420);
      gj_convolution3D_cp_element_group_421 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(421), clk => clk, reset => reset); --
    end block;
    -- CP-element group 422:  join  transition  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	418 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (1) 
      -- CP-element group 422: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(418) & convolution3D_CP_1120_elements(421);
      gj_convolution3D_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  merge  fork  transition  place  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	415 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423: 	425 
    -- CP-element group 423:  members (2) 
      -- CP-element group 423: 	 branch_block_stmt_436/merge_stmt_1559_PhiReqMerge
      -- CP-element group 423: 	 branch_block_stmt_436/merge_stmt_1559_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(423) <= OrReduce(convolution3D_CP_1120_elements(415) & convolution3D_CP_1120_elements(422));
    -- CP-element group 424:  transition  input  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	426 
    -- CP-element group 424:  members (1) 
      -- CP-element group 424: 	 branch_block_stmt_436/merge_stmt_1559_PhiAck/phi_stmt_1560_ack
      -- 
    phi_stmt_1560_ack_4222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1560_ack_0, ack => convolution3D_CP_1120_elements(424)); -- 
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	423 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (1) 
      -- CP-element group 425: 	 branch_block_stmt_436/merge_stmt_1559_PhiAck/phi_stmt_1567_ack
      -- 
    phi_stmt_1567_ack_4223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1567_ack_0, ack => convolution3D_CP_1120_elements(425)); -- 
    -- CP-element group 426:  join  fork  transition  place  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	424 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	317 
    -- CP-element group 426: 	322 
    -- CP-element group 426: 	323 
    -- CP-element group 426: 	324 
    -- CP-element group 426:  members (16) 
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_436/merge_stmt_1559__exit__
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616__entry__
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_update_start_
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_Update/$entry
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1610_Update/cr
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_Update/cr
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_Update/$entry
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/type_cast_1595_update_start_
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/RPIPE_maxpool_input_pipe_1588_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_436/assign_stmt_1580_to_assign_stmt_1616/$entry
      -- CP-element group 426: 	 branch_block_stmt_436/merge_stmt_1559_PhiAck/$exit
      -- 
    rr_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(426), ack => type_cast_1610_inst_req_0); -- 
    cr_3426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(426), ack => type_cast_1610_inst_req_1); -- 
    cr_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(426), ack => type_cast_1595_inst_req_1); -- 
    rr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(426), ack => RPIPE_maxpool_input_pipe_1588_inst_req_0); -- 
    convolution3D_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(424) & convolution3D_CP_1120_elements(425);
      gj_convolution3D_cp_element_group_426 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	327 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	429 
    -- CP-element group 427:  members (2) 
      -- CP-element group 427: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/$exit
      -- CP-element group 427: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Sample/ra
      -- 
    ra_4247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_0, ack => convolution3D_CP_1120_elements(427)); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	327 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (2) 
      -- CP-element group 428: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/$exit
      -- CP-element group 428: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/Update/ca
      -- 
    ca_4252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_1, ack => convolution3D_CP_1120_elements(428)); -- 
    -- CP-element group 429:  join  transition  place  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	427 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (8) 
      -- CP-element group 429: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/$exit
      -- CP-element group 429: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/$exit
      -- CP-element group 429: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/$exit
      -- CP-element group 429: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/$exit
      -- CP-element group 429: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_sources/type_cast_1627/SplitProtocol/$exit
      -- CP-element group 429: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1624/phi_stmt_1624_req
      -- CP-element group 429: 	 branch_block_stmt_436/merge_stmt_1623_PhiReqMerge
      -- CP-element group 429: 	 branch_block_stmt_436/merge_stmt_1623_PhiAck/$entry
      -- 
    phi_stmt_1624_req_4253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1624_req_4253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(429), ack => phi_stmt_1624_req_0); -- 
    convolution3D_cp_element_group_429: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_429"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(427) & convolution3D_CP_1120_elements(428);
      gj_convolution3D_cp_element_group_429 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(429), clk => clk, reset => reset); --
    end block;
    -- CP-element group 430:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	329 
    -- CP-element group 430: 	331 
    -- CP-element group 430: 	328 
    -- CP-element group 430: 	333 
    -- CP-element group 430:  members (29) 
      -- CP-element group 430: 	 branch_block_stmt_436/merge_stmt_1623__exit__
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662__entry__
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Update/word_access_complete/word_0/cr
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Update/word_access_complete/word_0/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_update_start_
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Update/word_access_complete/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/ptr_deref_1660_Update/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_complete/req
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_complete/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_Update/req
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_Update/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_Sample/req
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_final_index_sum_regn_update_start
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_scale_1/scale_rename_ack
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_scale_1/scale_rename_req
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_scale_1/$exit
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_scale_1/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_resize_1/index_resize_ack
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_resize_1/index_resize_req
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_resize_1/$exit
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_resize_1/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_computed_1
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_scaled_1
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/array_obj_ref_1656_index_resized_1
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1634_to_assign_stmt_1662/addr_of_1657_update_start_
      -- CP-element group 430: 	 branch_block_stmt_436/merge_stmt_1623_PhiAck/$exit
      -- CP-element group 430: 	 branch_block_stmt_436/merge_stmt_1623_PhiAck/phi_stmt_1624_ack
      -- 
    phi_stmt_1624_ack_4258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1624_ack_0, ack => convolution3D_CP_1120_elements(430)); -- 
    cr_3544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => ptr_deref_1660_store_0_req_1); -- 
    req_3494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => addr_of_1657_final_reg_req_1); -- 
    req_3479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => array_obj_ref_1656_index_offset_req_1); -- 
    req_3474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => array_obj_ref_1656_index_offset_req_0); -- 
    -- CP-element group 431:  merge  fork  transition  place  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	334 
    -- CP-element group 431: 	313 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	335 
    -- CP-element group 431: 	336 
    -- CP-element group 431:  members (13) 
      -- CP-element group 431: 	 branch_block_stmt_436/merge_stmt_1664__exit__
      -- CP-element group 431: 	 branch_block_stmt_436/call_stmt_1667__entry__
      -- CP-element group 431: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_sample_start_
      -- CP-element group 431: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_update_start_
      -- CP-element group 431: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_Sample/$entry
      -- CP-element group 431: 	 branch_block_stmt_436/call_stmt_1667/$entry
      -- CP-element group 431: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_Update/ccr
      -- CP-element group 431: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_Update/$entry
      -- CP-element group 431: 	 branch_block_stmt_436/call_stmt_1667/call_stmt_1667_Sample/crr
      -- CP-element group 431: 	 branch_block_stmt_436/merge_stmt_1664_PhiReqMerge
      -- CP-element group 431: 	 branch_block_stmt_436/merge_stmt_1664_PhiAck/$entry
      -- CP-element group 431: 	 branch_block_stmt_436/merge_stmt_1664_PhiAck/$exit
      -- CP-element group 431: 	 branch_block_stmt_436/merge_stmt_1664_PhiAck/dummy
      -- 
    ccr_3561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(431), ack => call_stmt_1667_call_req_1); -- 
    crr_3556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(431), ack => call_stmt_1667_call_req_0); -- 
    convolution3D_CP_1120_elements(431) <= OrReduce(convolution3D_CP_1120_elements(334) & convolution3D_CP_1120_elements(313));
    -- CP-element group 432:  transition  output  delay-element  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	349 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	436 
    -- CP-element group 432:  members (5) 
      -- CP-element group 432: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/$exit
      -- CP-element group 432: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1738/$exit
      -- CP-element group 432: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/$exit
      -- CP-element group 432: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1744_konst_delay_trans
      -- CP-element group 432: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_req
      -- 
    phi_stmt_1738_req_4280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1738_req_4280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(432), ack => phi_stmt_1738_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(432) is a control-delay.
    cp_element_432_delay: control_delay_element  generic map(name => " 432_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(349), ack => convolution3D_CP_1120_elements(432), clk => clk, reset =>reset);
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	361 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	435 
    -- CP-element group 433:  members (2) 
      -- CP-element group 433: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/Sample/$exit
      -- CP-element group 433: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/Sample/ra
      -- 
    ra_4300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1741_inst_ack_0, ack => convolution3D_CP_1120_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	361 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	435 
    -- CP-element group 434:  members (2) 
      -- CP-element group 434: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/Update/$exit
      -- CP-element group 434: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/Update/ca
      -- 
    ca_4305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1741_inst_ack_1, ack => convolution3D_CP_1120_elements(434)); -- 
    -- CP-element group 435:  join  transition  output  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	433 
    -- CP-element group 435: 	434 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (6) 
      -- CP-element group 435: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 435: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/$exit
      -- CP-element group 435: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/$exit
      -- CP-element group 435: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/$exit
      -- CP-element group 435: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_sources/type_cast_1741/SplitProtocol/$exit
      -- CP-element group 435: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1738/phi_stmt_1738_req
      -- 
    phi_stmt_1738_req_4306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1738_req_4306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(435), ack => phi_stmt_1738_req_0); -- 
    convolution3D_cp_element_group_435: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_435"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(433) & convolution3D_CP_1120_elements(434);
      gj_convolution3D_cp_element_group_435 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(435), clk => clk, reset => reset); --
    end block;
    -- CP-element group 436:  merge  transition  place  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	432 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436:  members (2) 
      -- CP-element group 436: 	 branch_block_stmt_436/merge_stmt_1737_PhiReqMerge
      -- CP-element group 436: 	 branch_block_stmt_436/merge_stmt_1737_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(436) <= OrReduce(convolution3D_CP_1120_elements(432) & convolution3D_CP_1120_elements(435));
    -- CP-element group 437:  fork  transition  place  input  output  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	356 
    -- CP-element group 437: 	357 
    -- CP-element group 437: 	358 
    -- CP-element group 437: 	350 
    -- CP-element group 437: 	351 
    -- CP-element group 437: 	352 
    -- CP-element group 437: 	353 
    -- CP-element group 437:  members (26) 
      -- CP-element group 437: 	 branch_block_stmt_436/merge_stmt_1737__exit__
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784__entry__
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_update_start_
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_Update/cr
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_Sample/rr
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_sample_start_
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/$entry
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_sample_start_
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_Update/$entry
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_update_start_
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_Sample/rr
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1758_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_Update/$entry
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/type_cast_1762_Update/cr
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_update_start_
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_Update/$entry
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1766_Update/ccr
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_sample_start_
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_update_start_
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_Sample/crr
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_Update/$entry
      -- CP-element group 437: 	 branch_block_stmt_436/assign_stmt_1750_to_assign_stmt_1784/call_stmt_1773_Update/ccr
      -- CP-element group 437: 	 branch_block_stmt_436/merge_stmt_1737_PhiAck/$exit
      -- CP-element group 437: 	 branch_block_stmt_436/merge_stmt_1737_PhiAck/phi_stmt_1738_ack
      -- 
    phi_stmt_1738_ack_4311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1738_ack_0, ack => convolution3D_CP_1120_elements(437)); -- 
    cr_3665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(437), ack => type_cast_1758_inst_req_1); -- 
    rr_3674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(437), ack => type_cast_1762_inst_req_0); -- 
    rr_3660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(437), ack => type_cast_1758_inst_req_0); -- 
    cr_3679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(437), ack => type_cast_1762_inst_req_1); -- 
    ccr_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(437), ack => call_stmt_1766_call_req_1); -- 
    crr_3702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(437), ack => call_stmt_1773_call_req_0); -- 
    ccr_3707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(437), ack => call_stmt_1773_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1014_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1208_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1510_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1134 : std_logic_vector(63 downto 0);
    signal R_indvar476_1308_resized : std_logic_vector(13 downto 0);
    signal R_indvar476_1308_scaled : std_logic_vector(13 downto 0);
    signal R_indvar490_812_resized : std_logic_vector(13 downto 0);
    signal R_indvar490_812_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1155_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1155_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1655_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1655_scaled : std_logic_vector(13 downto 0);
    signal add117_661 : std_logic_vector(15 downto 0);
    signal add135_692 : std_logic_vector(15 downto 0);
    signal add1519x_xi434_1640 : std_logic_vector(63 downto 0);
    signal add1519x_xi_1140 : std_logic_vector(63 downto 0);
    signal add166_846 : std_logic_vector(63 downto 0);
    signal add176_867 : std_logic_vector(63 downto 0);
    signal add186_888 : std_logic_vector(63 downto 0);
    signal add196_909 : std_logic_vector(63 downto 0);
    signal add206_930 : std_logic_vector(63 downto 0);
    signal add216_951 : std_logic_vector(63 downto 0);
    signal add226_972 : std_logic_vector(63 downto 0);
    signal add273_1342 : std_logic_vector(63 downto 0);
    signal add27_506 : std_logic_vector(15 downto 0);
    signal add283_1363 : std_logic_vector(63 downto 0);
    signal add293_1384 : std_logic_vector(63 downto 0);
    signal add303_1405 : std_logic_vector(63 downto 0);
    signal add313_1426 : std_logic_vector(63 downto 0);
    signal add323_1447 : std_logic_vector(63 downto 0);
    signal add333_1468 : std_logic_vector(63 downto 0);
    signal add45_537 : std_logic_vector(15 downto 0);
    signal add63_568 : std_logic_vector(15 downto 0);
    signal add81_599 : std_logic_vector(15 downto 0);
    signal add99_630 : std_logic_vector(15 downto 0);
    signal add_475 : std_logic_vector(31 downto 0);
    signal addx_xi425_1601 : std_logic_vector(63 downto 0);
    signal addx_xi_1101 : std_logic_vector(63 downto 0);
    signal and343_1528 : std_logic_vector(63 downto 0);
    signal and_1032 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1156_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1156_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1156_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1156_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1156_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1156_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1656_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1656_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1656_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1656_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1656_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1656_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_813_root_address : std_logic_vector(13 downto 0);
    signal arrayidx237_1158 : std_logic_vector(31 downto 0);
    signal arrayidx337_1311 : std_logic_vector(31 downto 0);
    signal arrayidx352_1658 : std_logic_vector(31 downto 0);
    signal arrayidx_815 : std_logic_vector(31 downto 0);
    signal call104_633 : std_logic_vector(7 downto 0);
    signal call113_649 : std_logic_vector(7 downto 0);
    signal call122_664 : std_logic_vector(7 downto 0);
    signal call131_680 : std_logic_vector(7 downto 0);
    signal call14_478 : std_logic_vector(7 downto 0);
    signal call153_818 : std_logic_vector(7 downto 0);
    signal call161_834 : std_logic_vector(7 downto 0);
    signal call171_855 : std_logic_vector(7 downto 0);
    signal call181_876 : std_logic_vector(7 downto 0);
    signal call191_897 : std_logic_vector(7 downto 0);
    signal call201_918 : std_logic_vector(7 downto 0);
    signal call211_939 : std_logic_vector(7 downto 0);
    signal call221_960 : std_logic_vector(7 downto 0);
    signal call23_494 : std_logic_vector(7 downto 0);
    signal call260_1314 : std_logic_vector(7 downto 0);
    signal call268_1330 : std_logic_vector(7 downto 0);
    signal call278_1351 : std_logic_vector(7 downto 0);
    signal call288_1372 : std_logic_vector(7 downto 0);
    signal call298_1393 : std_logic_vector(7 downto 0);
    signal call308_1414 : std_logic_vector(7 downto 0);
    signal call318_1435 : std_logic_vector(7 downto 0);
    signal call328_1456 : std_logic_vector(7 downto 0);
    signal call32_509 : std_logic_vector(7 downto 0);
    signal call355_1667 : std_logic_vector(63 downto 0);
    signal call410_1799 : std_logic_vector(63 downto 0);
    signal call41_525 : std_logic_vector(7 downto 0);
    signal call50_540 : std_logic_vector(7 downto 0);
    signal call59_556 : std_logic_vector(7 downto 0);
    signal call68_571 : std_logic_vector(7 downto 0);
    signal call6_463 : std_logic_vector(7 downto 0);
    signal call77_587 : std_logic_vector(7 downto 0);
    signal call86_602 : std_logic_vector(7 downto 0);
    signal call95_618 : std_logic_vector(7 downto 0);
    signal call_447 : std_logic_vector(7 downto 0);
    signal callx_xi423_1589 : std_logic_vector(7 downto 0);
    signal callx_xi_1089 : std_logic_vector(7 downto 0);
    signal cmp255443_1216 : std_logic_vector(0 downto 0);
    signal cmp447_722 : std_logic_vector(0 downto 0);
    signal cmpx_xi428_1616 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1116 : std_logic_vector(0 downto 0);
    signal conv109_640 : std_logic_vector(15 downto 0);
    signal conv116_656 : std_logic_vector(15 downto 0);
    signal conv127_671 : std_logic_vector(15 downto 0);
    signal conv134_687 : std_logic_vector(15 downto 0);
    signal conv141_696 : std_logic_vector(31 downto 0);
    signal conv143_700 : std_logic_vector(31 downto 0);
    signal conv145_716 : std_logic_vector(63 downto 0);
    signal conv156_825 : std_logic_vector(63 downto 0);
    signal conv165_841 : std_logic_vector(63 downto 0);
    signal conv175_862 : std_logic_vector(63 downto 0);
    signal conv185_883 : std_logic_vector(63 downto 0);
    signal conv195_904 : std_logic_vector(63 downto 0);
    signal conv19_485 : std_logic_vector(15 downto 0);
    signal conv205_925 : std_logic_vector(63 downto 0);
    signal conv215_946 : std_logic_vector(63 downto 0);
    signal conv225_967 : std_logic_vector(63 downto 0);
    signal conv239_1168 : std_logic_vector(63 downto 0);
    signal conv241_1172 : std_logic_vector(63 downto 0);
    signal conv244_1176 : std_logic_vector(63 downto 0);
    signal conv247_1180 : std_logic_vector(63 downto 0);
    signal conv249_1210 : std_logic_vector(63 downto 0);
    signal conv263_1321 : std_logic_vector(63 downto 0);
    signal conv26_501 : std_logic_vector(15 downto 0);
    signal conv272_1337 : std_logic_vector(63 downto 0);
    signal conv282_1358 : std_logic_vector(63 downto 0);
    signal conv292_1379 : std_logic_vector(63 downto 0);
    signal conv2x_xi418_1551 : std_logic_vector(31 downto 0);
    signal conv2x_xi_1051 : std_logic_vector(31 downto 0);
    signal conv302_1400 : std_logic_vector(63 downto 0);
    signal conv312_1421 : std_logic_vector(63 downto 0);
    signal conv322_1442 : std_logic_vector(63 downto 0);
    signal conv332_1463 : std_logic_vector(63 downto 0);
    signal conv356_1796 : std_logic_vector(63 downto 0);
    signal conv37_516 : std_logic_vector(15 downto 0);
    signal conv381_1759 : std_logic_vector(63 downto 0);
    signal conv387_1763 : std_logic_vector(63 downto 0);
    signal conv3_454 : std_logic_vector(31 downto 0);
    signal conv411_1804 : std_logic_vector(63 downto 0);
    signal conv44_532 : std_logic_vector(15 downto 0);
    signal conv55_547 : std_logic_vector(15 downto 0);
    signal conv62_563 : std_logic_vector(15 downto 0);
    signal conv73_578 : std_logic_vector(15 downto 0);
    signal conv80_594 : std_logic_vector(15 downto 0);
    signal conv8x_xi424_1596 : std_logic_vector(63 downto 0);
    signal conv8x_xi_1096 : std_logic_vector(63 downto 0);
    signal conv91_609 : std_logic_vector(15 downto 0);
    signal conv98_625 : std_logic_vector(15 downto 0);
    signal conv9_470 : std_logic_vector(31 downto 0);
    signal convx_xi427_1611 : std_logic_vector(31 downto 0);
    signal convx_xi_1111 : std_logic_vector(31 downto 0);
    signal elementx_x024x_xi422_1567 : std_logic_vector(63 downto 0);
    signal elementx_x024x_xi_1067 : std_logic_vector(63 downto 0);
    signal exitcond32_987 : std_logic_vector(0 downto 0);
    signal exitcond5_1784 : std_logic_vector(0 downto 0);
    signal exitcond_1483 : std_logic_vector(0 downto 0);
    signal iNsTr_126_1547 : std_logic_vector(63 downto 0);
    signal iNsTr_134_1586 : std_logic_vector(15 downto 0);
    signal iNsTr_144_1634 : std_logic_vector(63 downto 0);
    signal iNsTr_86_1086 : std_logic_vector(15 downto 0);
    signal indvar476_1297 : std_logic_vector(63 downto 0);
    signal indvar490_801 : std_logic_vector(63 downto 0);
    signal indvar_1738 : std_logic_vector(31 downto 0);
    signal indvarx_xnext477_1478 : std_logic_vector(63 downto 0);
    signal indvarx_xnext491_982 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1779 : std_logic_vector(31 downto 0);
    signal ix_x0x_xlcssa_1019 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1515 : std_logic_vector(63 downto 0);
    signal mul144_710 : std_logic_vector(31 downto 0);
    signal mul242_1185 : std_logic_vector(63 downto 0);
    signal mul245_1190 : std_logic_vector(63 downto 0);
    signal mul248_1195 : std_logic_vector(63 downto 0);
    signal mul362_1673 : std_logic_vector(15 downto 0);
    signal mul375_1678 : std_logic_vector(15 downto 0);
    signal mul380_1750 : std_logic_vector(31 downto 0);
    signal mul386_1755 : std_logic_vector(31 downto 0);
    signal mul_705 : std_logic_vector(31 downto 0);
    signal nx_x025x_xi421_1560 : std_logic_vector(15 downto 0);
    signal nx_x025x_xi_1060 : std_logic_vector(15 downto 0);
    signal phitmp451_1512 : std_logic_vector(63 downto 0);
    signal phitmp_1016 : std_logic_vector(63 downto 0);
    signal ptr_deref_1160_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1160_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1160_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1470_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1470_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1470_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1470_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1470_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1470_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1660_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1660_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1660_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1660_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1660_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1660_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_974_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_974_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_974_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_974_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_974_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_974_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_1201 : std_logic_vector(63 downto 0);
    signal sh_promx_xi435_1646 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1146 : std_logic_vector(63 downto 0);
    signal shl110_646 : std_logic_vector(15 downto 0);
    signal shl11x_xi426_1607 : std_logic_vector(63 downto 0);
    signal shl11x_xi426x_xlcssa_1624 : std_logic_vector(63 downto 0);
    signal shl11x_xi_1107 : std_logic_vector(63 downto 0);
    signal shl11x_xix_xlcssa_1124 : std_logic_vector(63 downto 0);
    signal shl128_677 : std_logic_vector(15 downto 0);
    signal shl158_831 : std_logic_vector(63 downto 0);
    signal shl168_852 : std_logic_vector(63 downto 0);
    signal shl178_873 : std_logic_vector(63 downto 0);
    signal shl17x_xi436_1651 : std_logic_vector(63 downto 0);
    signal shl17x_xi_1151 : std_logic_vector(63 downto 0);
    signal shl188_894 : std_logic_vector(63 downto 0);
    signal shl198_915 : std_logic_vector(63 downto 0);
    signal shl208_936 : std_logic_vector(63 downto 0);
    signal shl20_491 : std_logic_vector(15 downto 0);
    signal shl218_957 : std_logic_vector(63 downto 0);
    signal shl265_1327 : std_logic_vector(63 downto 0);
    signal shl275_1348 : std_logic_vector(63 downto 0);
    signal shl285_1369 : std_logic_vector(63 downto 0);
    signal shl295_1390 : std_logic_vector(63 downto 0);
    signal shl305_1411 : std_logic_vector(63 downto 0);
    signal shl315_1432 : std_logic_vector(63 downto 0);
    signal shl325_1453 : std_logic_vector(63 downto 0);
    signal shl38_522 : std_logic_vector(15 downto 0);
    signal shl56_553 : std_logic_vector(15 downto 0);
    signal shl74_584 : std_logic_vector(15 downto 0);
    signal shl92_615 : std_logic_vector(15 downto 0);
    signal shl_460 : std_logic_vector(31 downto 0);
    signal shlx_xi419_1557 : std_logic_vector(31 downto 0);
    signal shlx_xi_1057 : std_logic_vector(31 downto 0);
    signal sub395_1701 : std_logic_vector(15 downto 0);
    signal sub415_1809 : std_logic_vector(63 downto 0);
    signal sub_1695 : std_logic_vector(15 downto 0);
    signal tmp12_1239 : std_logic_vector(63 downto 0);
    signal tmp13_1243 : std_logic_vector(63 downto 0);
    signal tmp14_1248 : std_logic_vector(63 downto 0);
    signal tmp15_1252 : std_logic_vector(63 downto 0);
    signal tmp16_1257 : std_logic_vector(63 downto 0);
    signal tmp17_1261 : std_logic_vector(63 downto 0);
    signal tmp18_1266 : std_logic_vector(63 downto 0);
    signal tmp19_1270 : std_logic_vector(31 downto 0);
    signal tmp20_1275 : std_logic_vector(63 downto 0);
    signal tmp21_1281 : std_logic_vector(63 downto 0);
    signal tmp22_1287 : std_logic_vector(0 downto 0);
    signal tmp24_760 : std_logic_vector(31 downto 0);
    signal tmp25_765 : std_logic_vector(31 downto 0);
    signal tmp26_769 : std_logic_vector(31 downto 0);
    signal tmp27_774 : std_logic_vector(31 downto 0);
    signal tmp28_779 : std_logic_vector(63 downto 0);
    signal tmp29_785 : std_logic_vector(63 downto 0);
    signal tmp30_791 : std_logic_vector(0 downto 0);
    signal tmp3_1711 : std_logic_vector(31 downto 0);
    signal tmp452_1580 : std_logic_vector(15 downto 0);
    signal tmp453_1707 : std_logic_vector(15 downto 0);
    signal tmp471_1229 : std_logic_vector(63 downto 0);
    signal tmp472_1235 : std_logic_vector(0 downto 0);
    signal tmp473_1503 : std_logic_vector(63 downto 0);
    signal tmp480_734 : std_logic_vector(31 downto 0);
    signal tmp482_739 : std_logic_vector(31 downto 0);
    signal tmp483_744 : std_logic_vector(63 downto 0);
    signal tmp484_750 : std_logic_vector(63 downto 0);
    signal tmp485_756 : std_logic_vector(0 downto 0);
    signal tmp487_1007 : std_logic_vector(63 downto 0);
    signal tmp4_1717 : std_logic_vector(31 downto 0);
    signal tmp6_1721 : std_logic_vector(31 downto 0);
    signal tmp7_1726 : std_logic_vector(15 downto 0);
    signal tmp8_1730 : std_logic_vector(31 downto 0);
    signal tmp9_1735 : std_logic_vector(31 downto 0);
    signal tmp_1080 : std_logic_vector(15 downto 0);
    signal tobool344_1534 : std_logic_vector(0 downto 0);
    signal tobool_1038 : std_logic_vector(0 downto 0);
    signal type_cast_1005_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1010_wire : std_logic_vector(63 downto 0);
    signal type_cast_1013_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1022_wire : std_logic_vector(63 downto 0);
    signal type_cast_1025_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1030_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1036_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1049_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1055_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1064_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1066_wire : std_logic_vector(15 downto 0);
    signal type_cast_1071_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1073_wire : std_logic_vector(63 downto 0);
    signal type_cast_1078_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1084_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1105_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1127_wire : std_logic_vector(63 downto 0);
    signal type_cast_1132_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1138_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1199_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1204_wire : std_logic_vector(63 downto 0);
    signal type_cast_1207_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1214_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1227_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1233_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1273_wire : std_logic_vector(63 downto 0);
    signal type_cast_1279_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1285_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1292_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1301_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1303_wire : std_logic_vector(63 downto 0);
    signal type_cast_1325_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1346_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1367_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1388_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1409_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1430_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1451_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1476_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1495_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1501_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1506_wire : std_logic_vector(63 downto 0);
    signal type_cast_1509_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1519_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1521_wire : std_logic_vector(63 downto 0);
    signal type_cast_1526_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1532_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1545_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1555_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1564_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1566_wire : std_logic_vector(15 downto 0);
    signal type_cast_1571_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1573_wire : std_logic_vector(63 downto 0);
    signal type_cast_1578_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1584_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1605_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1627_wire : std_logic_vector(63 downto 0);
    signal type_cast_1632_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1638_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1644_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1684_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1688_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1693_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1699_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1705_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1715_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1741_wire : std_logic_vector(31 downto 0);
    signal type_cast_1744_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1777_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1794_wire : std_logic_vector(63 downto 0);
    signal type_cast_1802_wire : std_logic_vector(63 downto 0);
    signal type_cast_439_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_443_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_458_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_489_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_551_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_613_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_644_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_675_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_714_wire : std_logic_vector(63 downto 0);
    signal type_cast_720_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_742_wire : std_logic_vector(63 downto 0);
    signal type_cast_748_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_754_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_777_wire : std_logic_vector(63 downto 0);
    signal type_cast_783_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_789_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_805_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_807_wire : std_logic_vector(63 downto 0);
    signal type_cast_829_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_850_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_871_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_913_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_934_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_955_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_980_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_999_wire_constant : std_logic_vector(63 downto 0);
    signal umax23_1294 : std_logic_vector(63 downto 0);
    signal umax31_798 : std_logic_vector(63 downto 0);
    signal umax486_1001 : std_logic_vector(63 downto 0);
    signal umax_1497 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1156_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1156_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1156_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1156_resized_base_address <= "00000000000000";
    array_obj_ref_1309_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1309_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1309_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1309_resized_base_address <= "00000000000000";
    array_obj_ref_1656_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1656_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1656_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1656_resized_base_address <= "00000000000000";
    array_obj_ref_813_constant_part_of_offset <= "00000000000000";
    array_obj_ref_813_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_813_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_813_resized_base_address <= "00000000000000";
    ptr_deref_1160_word_offset_0 <= "00000000000000";
    ptr_deref_1470_word_offset_0 <= "00000000000000";
    ptr_deref_1660_word_offset_0 <= "00000000000000";
    ptr_deref_974_word_offset_0 <= "00000000000000";
    type_cast_1005_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1013_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1025_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1030_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1036_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1049_wire_constant <= "00000000000000000000000000000001";
    type_cast_1055_wire_constant <= "00000000000000000000000000000110";
    type_cast_1064_wire_constant <= "0000000000000000";
    type_cast_1071_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1078_wire_constant <= "0000000000000001";
    type_cast_1084_wire_constant <= "0000000000000001";
    type_cast_1105_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1132_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1138_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1144_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1199_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1207_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1214_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1227_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1233_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1279_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1285_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1292_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1301_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1325_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1346_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1367_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1388_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1409_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1430_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1451_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1476_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1495_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1501_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1509_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1519_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1526_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1532_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1545_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1555_wire_constant <= "00000000000000000000000000000110";
    type_cast_1564_wire_constant <= "0000000000000000";
    type_cast_1571_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1578_wire_constant <= "0000000000000001";
    type_cast_1584_wire_constant <= "0000000000000001";
    type_cast_1605_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1632_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1638_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1644_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1684_wire_constant <= "11001000";
    type_cast_1688_wire_constant <= "11001000";
    type_cast_1693_wire_constant <= "1111111111111111";
    type_cast_1699_wire_constant <= "1111111111111111";
    type_cast_1705_wire_constant <= "1111111111111111";
    type_cast_1715_wire_constant <= "00000000000000000000000000000001";
    type_cast_1744_wire_constant <= "00000000000000000000000000000000";
    type_cast_1777_wire_constant <= "00000000000000000000000000000001";
    type_cast_439_wire_constant <= "01100100";
    type_cast_443_wire_constant <= "01100100";
    type_cast_458_wire_constant <= "00000000000000000000000000001000";
    type_cast_489_wire_constant <= "0000000000001000";
    type_cast_520_wire_constant <= "0000000000001000";
    type_cast_551_wire_constant <= "0000000000001000";
    type_cast_582_wire_constant <= "0000000000001000";
    type_cast_613_wire_constant <= "0000000000001000";
    type_cast_644_wire_constant <= "0000000000001000";
    type_cast_675_wire_constant <= "0000000000001000";
    type_cast_720_wire_constant <= "00000000000000000000000000000011";
    type_cast_748_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_754_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_783_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_789_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_796_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_805_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_829_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_850_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_871_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_892_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_913_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_934_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_955_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_980_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_999_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1019: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1022_wire & type_cast_1025_wire_constant;
      req <= phi_stmt_1019_req_0 & phi_stmt_1019_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1019",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1019_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_1019,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1019
    phi_stmt_1060: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1064_wire_constant & type_cast_1066_wire;
      req <= phi_stmt_1060_req_0 & phi_stmt_1060_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1060",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1060_ack_0,
          idata => idata,
          odata => nx_x025x_xi_1060,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1060
    phi_stmt_1067: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1071_wire_constant & type_cast_1073_wire;
      req <= phi_stmt_1067_req_0 & phi_stmt_1067_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1067",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1067_ack_0,
          idata => idata,
          odata => elementx_x024x_xi_1067,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1067
    phi_stmt_1124: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1127_wire;
      req(0) <= phi_stmt_1124_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1124",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1124_ack_0,
          idata => idata,
          odata => shl11x_xix_xlcssa_1124,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1124
    phi_stmt_1297: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1301_wire_constant & type_cast_1303_wire;
      req <= phi_stmt_1297_req_0 & phi_stmt_1297_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1297",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1297_ack_0,
          idata => idata,
          odata => indvar476_1297,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1297
    phi_stmt_1515: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1519_wire_constant & type_cast_1521_wire;
      req <= phi_stmt_1515_req_0 & phi_stmt_1515_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1515",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1515_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1515,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1515
    phi_stmt_1560: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1564_wire_constant & type_cast_1566_wire;
      req <= phi_stmt_1560_req_0 & phi_stmt_1560_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1560",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1560_ack_0,
          idata => idata,
          odata => nx_x025x_xi421_1560,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1560
    phi_stmt_1567: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1571_wire_constant & type_cast_1573_wire;
      req <= phi_stmt_1567_req_0 & phi_stmt_1567_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1567",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1567_ack_0,
          idata => idata,
          odata => elementx_x024x_xi422_1567,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1567
    phi_stmt_1624: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1627_wire;
      req(0) <= phi_stmt_1624_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1624",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1624_ack_0,
          idata => idata,
          odata => shl11x_xi426x_xlcssa_1624,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1624
    phi_stmt_1738: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1741_wire & type_cast_1744_wire_constant;
      req <= phi_stmt_1738_req_0 & phi_stmt_1738_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1738",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1738_ack_0,
          idata => idata,
          odata => indvar_1738,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1738
    phi_stmt_801: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_805_wire_constant & type_cast_807_wire;
      req <= phi_stmt_801_req_0 & phi_stmt_801_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_801",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_801_ack_0,
          idata => idata,
          odata => indvar490_801,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_801
    -- flow-through select operator MUX_1000_inst
    umax486_1001 <= tmp484_750 when (tmp485_756(0) /=  '0') else type_cast_999_wire_constant;
    -- flow-through select operator MUX_1293_inst
    umax23_1294 <= tmp21_1281 when (tmp22_1287(0) /=  '0') else type_cast_1292_wire_constant;
    -- flow-through select operator MUX_1496_inst
    umax_1497 <= tmp471_1229 when (tmp472_1235(0) /=  '0') else type_cast_1495_wire_constant;
    -- flow-through select operator MUX_797_inst
    umax31_798 <= tmp29_785 when (tmp30_791(0) /=  '0') else type_cast_796_wire_constant;
    addr_of_1157_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1157_final_reg_req_0;
      addr_of_1157_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1157_final_reg_req_1;
      addr_of_1157_final_reg_ack_1<= rack(0);
      addr_of_1157_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1157_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1156_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx237_1158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1310_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1310_final_reg_req_0;
      addr_of_1310_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1310_final_reg_req_1;
      addr_of_1310_final_reg_ack_1<= rack(0);
      addr_of_1310_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1310_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1309_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx337_1311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1657_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1657_final_reg_req_0;
      addr_of_1657_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1657_final_reg_req_1;
      addr_of_1657_final_reg_ack_1<= rack(0);
      addr_of_1657_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1657_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1656_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx352_1658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_814_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_814_final_reg_req_0;
      addr_of_814_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_814_final_reg_req_1;
      addr_of_814_final_reg_ack_1<= rack(0);
      addr_of_814_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_814_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_813_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1010_inst
    process(tmp487_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp487_1007(63 downto 0);
      type_cast_1010_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1015_inst
    process(ASHR_i64_i64_1014_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1014_wire(63 downto 0);
      phitmp_1016 <= tmp_var; -- 
    end process;
    type_cast_1022_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1022_inst_req_0;
      type_cast_1022_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1022_inst_req_1;
      type_cast_1022_inst_ack_1<= rack(0);
      type_cast_1022_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1022_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_1016,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1022_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1066_inst_req_0;
      type_cast_1066_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1066_inst_req_1;
      type_cast_1066_inst_ack_1<= rack(0);
      type_cast_1066_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1066_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_86_1086,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1066_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1073_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1073_inst_req_0;
      type_cast_1073_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1073_inst_req_1;
      type_cast_1073_inst_ack_1<= rack(0);
      type_cast_1073_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1073_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl11x_xi_1107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1073_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1095_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1095_inst_req_0;
      type_cast_1095_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1095_inst_req_1;
      type_cast_1095_inst_ack_1<= rack(0);
      type_cast_1095_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1095_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1089,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8x_xi_1096,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1110_inst_req_0;
      type_cast_1110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1110_inst_req_1;
      type_cast_1110_inst_ack_1<= rack(0);
      type_cast_1110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1080,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1127_inst_req_0;
      type_cast_1127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1127_inst_req_1;
      type_cast_1127_inst_ack_1<= rack(0);
      type_cast_1127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl11x_xi_1107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1127_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1167_inst_req_0;
      type_cast_1167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1167_inst_req_1;
      type_cast_1167_inst_ack_1<= rack(0);
      type_cast_1167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add45_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv239_1168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1171_inst_req_0;
      type_cast_1171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1171_inst_req_1;
      type_cast_1171_inst_ack_1<= rack(0);
      type_cast_1171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1171_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_1172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1175_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1175_inst_req_0;
      type_cast_1175_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1175_inst_req_1;
      type_cast_1175_inst_ack_1<= rack(0);
      type_cast_1175_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1175_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv244_1176,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1179_inst_req_0;
      type_cast_1179_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1179_inst_req_1;
      type_cast_1179_inst_ack_1<= rack(0);
      type_cast_1179_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1179_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add99_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv247_1180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1204_inst
    process(sext_1201) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1201(63 downto 0);
      type_cast_1204_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1209_inst
    process(ASHR_i64_i64_1208_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1208_wire(63 downto 0);
      conv249_1210 <= tmp_var; -- 
    end process;
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add99_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1242_inst_req_0;
      type_cast_1242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1242_inst_req_1;
      type_cast_1242_inst_ack_1<= rack(0);
      type_cast_1242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1242_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add45_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1251_inst_req_0;
      type_cast_1251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1251_inst_req_1;
      type_cast_1251_inst_ack_1<= rack(0);
      type_cast_1251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_1252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1260_inst_req_0;
      type_cast_1260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1260_inst_req_1;
      type_cast_1260_inst_ack_1<= rack(0);
      type_cast_1260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp17_1261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1269_inst_req_0;
      type_cast_1269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1269_inst_req_1;
      type_cast_1269_inst_ack_1<= rack(0);
      type_cast_1269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp18_1266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp19_1270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1274_inst_req_0;
      type_cast_1274_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1274_inst_req_1;
      type_cast_1274_inst_ack_1<= rack(0);
      type_cast_1274_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1274_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1273_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1275,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1303_inst_req_0;
      type_cast_1303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1303_inst_req_1;
      type_cast_1303_inst_ack_1<= rack(0);
      type_cast_1303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext477_1478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1303_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1320_inst_req_0;
      type_cast_1320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1320_inst_req_1;
      type_cast_1320_inst_ack_1<= rack(0);
      type_cast_1320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call260_1314,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv263_1321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1336_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1336_inst_req_0;
      type_cast_1336_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1336_inst_req_1;
      type_cast_1336_inst_ack_1<= rack(0);
      type_cast_1336_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1336_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call268_1330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv272_1337,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1357_inst_req_0;
      type_cast_1357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1357_inst_req_1;
      type_cast_1357_inst_ack_1<= rack(0);
      type_cast_1357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call278_1351,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv282_1358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1378_inst_req_0;
      type_cast_1378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1378_inst_req_1;
      type_cast_1378_inst_ack_1<= rack(0);
      type_cast_1378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call288_1372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv292_1379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1399_inst_req_0;
      type_cast_1399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1399_inst_req_1;
      type_cast_1399_inst_ack_1<= rack(0);
      type_cast_1399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1399_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call298_1393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv302_1400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1420_inst_req_0;
      type_cast_1420_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1420_inst_req_1;
      type_cast_1420_inst_ack_1<= rack(0);
      type_cast_1420_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1420_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call308_1414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv312_1421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1441_inst_req_0;
      type_cast_1441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1441_inst_req_1;
      type_cast_1441_inst_ack_1<= rack(0);
      type_cast_1441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call318_1435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1462_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1462_inst_req_0;
      type_cast_1462_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1462_inst_req_1;
      type_cast_1462_inst_ack_1<= rack(0);
      type_cast_1462_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1462_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call328_1456,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv332_1463,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1506_inst
    process(tmp473_1503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp473_1503(63 downto 0);
      type_cast_1506_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1511_inst
    process(ASHR_i64_i64_1510_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1510_wire(63 downto 0);
      phitmp451_1512 <= tmp_var; -- 
    end process;
    type_cast_1521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1521_inst_req_0;
      type_cast_1521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1521_inst_req_1;
      type_cast_1521_inst_ack_1<= rack(0);
      type_cast_1521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp451_1512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1521_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1550_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1550_inst_req_0;
      type_cast_1550_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1550_inst_req_1;
      type_cast_1550_inst_ack_1<= rack(0);
      type_cast_1550_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1550_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_126_1547,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi418_1551,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1566_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1566_inst_req_0;
      type_cast_1566_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1566_inst_req_1;
      type_cast_1566_inst_ack_1<= rack(0);
      type_cast_1566_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1566_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_134_1586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1566_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1573_inst_req_0;
      type_cast_1573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1573_inst_req_1;
      type_cast_1573_inst_ack_1<= rack(0);
      type_cast_1573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl11x_xi426_1607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1573_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1595_inst_req_0;
      type_cast_1595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1595_inst_req_1;
      type_cast_1595_inst_ack_1<= rack(0);
      type_cast_1595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi423_1589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8x_xi424_1596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1610_inst_req_0;
      type_cast_1610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1610_inst_req_1;
      type_cast_1610_inst_ack_1<= rack(0);
      type_cast_1610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp452_1580,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi427_1611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1627_inst_req_0;
      type_cast_1627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1627_inst_req_1;
      type_cast_1627_inst_ack_1<= rack(0);
      type_cast_1627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl11x_xi426_1607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1627_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1710_inst_req_0;
      type_cast_1710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1710_inst_req_1;
      type_cast_1710_inst_ack_1<= rack(0);
      type_cast_1710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp453_1707,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1720_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1720_inst_req_0;
      type_cast_1720_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1720_inst_req_1;
      type_cast_1720_inst_ack_1<= rack(0);
      type_cast_1720_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1720_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_1721,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1729_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1729_inst_req_0;
      type_cast_1729_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1729_inst_req_1;
      type_cast_1729_inst_ack_1<= rack(0);
      type_cast_1729_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1729_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_1726,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_1730,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1741_inst_req_0;
      type_cast_1741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1741_inst_req_1;
      type_cast_1741_inst_ack_1<= rack(0);
      type_cast_1741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1741_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1758_inst_req_0;
      type_cast_1758_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1758_inst_req_1;
      type_cast_1758_inst_ack_1<= rack(0);
      type_cast_1758_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1758_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul380_1750,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv381_1759,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1762_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1762_inst_req_0;
      type_cast_1762_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1762_inst_req_1;
      type_cast_1762_inst_ack_1<= rack(0);
      type_cast_1762_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1762_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul386_1755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv387_1763,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1795_inst_req_0;
      type_cast_1795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1795_inst_req_1;
      type_cast_1795_inst_ack_1<= rack(0);
      type_cast_1795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1794_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv356_1796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1803_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1803_inst_req_0;
      type_cast_1803_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1803_inst_req_1;
      type_cast_1803_inst_ack_1<= rack(0);
      type_cast_1803_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1803_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1802_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv411_1804,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_453_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_453_inst_req_0;
      type_cast_453_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_453_inst_req_1;
      type_cast_453_inst_ack_1<= rack(0);
      type_cast_453_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_453_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_447,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_454,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_469_inst_req_0;
      type_cast_469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_469_inst_req_1;
      type_cast_469_inst_ack_1<= rack(0);
      type_cast_469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_484_inst_req_0;
      type_cast_484_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_484_inst_req_1;
      type_cast_484_inst_ack_1<= rack(0);
      type_cast_484_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_484_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_485,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_500_inst_req_0;
      type_cast_500_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_500_inst_req_1;
      type_cast_500_inst_ack_1<= rack(0);
      type_cast_500_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_500_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_501,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_515_inst_req_0;
      type_cast_515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_515_inst_req_1;
      type_cast_515_inst_ack_1<= rack(0);
      type_cast_515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_509,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_531_inst_req_0;
      type_cast_531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_531_inst_req_1;
      type_cast_531_inst_ack_1<= rack(0);
      type_cast_531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_546_inst_req_0;
      type_cast_546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_546_inst_req_1;
      type_cast_546_inst_ack_1<= rack(0);
      type_cast_546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_546_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_540,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv55_547,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_562_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_562_inst_req_0;
      type_cast_562_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_562_inst_req_1;
      type_cast_562_inst_ack_1<= rack(0);
      type_cast_562_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_562_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call59_556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_563,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_577_inst_req_0;
      type_cast_577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_577_inst_req_1;
      type_cast_577_inst_ack_1<= rack(0);
      type_cast_577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_593_inst_req_0;
      type_cast_593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_593_inst_req_1;
      type_cast_593_inst_ack_1<= rack(0);
      type_cast_593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call77_587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_608_inst_req_0;
      type_cast_608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_608_inst_req_1;
      type_cast_608_inst_ack_1<= rack(0);
      type_cast_608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call86_602,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_609,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_624_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_624_inst_req_0;
      type_cast_624_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_624_inst_req_1;
      type_cast_624_inst_ack_1<= rack(0);
      type_cast_624_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_624_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_625,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_639_inst_req_0;
      type_cast_639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_639_inst_req_1;
      type_cast_639_inst_ack_1<= rack(0);
      type_cast_639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call104_633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_655_inst_req_0;
      type_cast_655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_655_inst_req_1;
      type_cast_655_inst_ack_1<= rack(0);
      type_cast_655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call113_649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_656,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_670_inst_req_0;
      type_cast_670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_670_inst_req_1;
      type_cast_670_inst_ack_1<= rack(0);
      type_cast_670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call122_664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_686_inst_req_0;
      type_cast_686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_686_inst_req_1;
      type_cast_686_inst_ack_1<= rack(0);
      type_cast_686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call131_680,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_695_inst_req_0;
      type_cast_695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_695_inst_req_1;
      type_cast_695_inst_ack_1<= rack(0);
      type_cast_695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add27_506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_699_inst_req_0;
      type_cast_699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_699_inst_req_1;
      type_cast_699_inst_ack_1<= rack(0);
      type_cast_699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add45_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_715_inst_req_0;
      type_cast_715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_715_inst_req_1;
      type_cast_715_inst_ack_1<= rack(0);
      type_cast_715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_714_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_743_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_743_inst_req_0;
      type_cast_743_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_743_inst_req_1;
      type_cast_743_inst_ack_1<= rack(0);
      type_cast_743_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_743_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_742_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp483_744,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_759_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_759_inst_req_0;
      type_cast_759_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_759_inst_req_1;
      type_cast_759_inst_ack_1<= rack(0);
      type_cast_759_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_759_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add27_506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_760,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_768_inst_req_0;
      type_cast_768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_768_inst_req_1;
      type_cast_768_inst_ack_1<= rack(0);
      type_cast_768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add45_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp26_769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_778_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_778_inst_req_0;
      type_cast_778_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_778_inst_req_1;
      type_cast_778_inst_ack_1<= rack(0);
      type_cast_778_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_778_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_777_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp28_779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_807_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_807_inst_req_0;
      type_cast_807_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_807_inst_req_1;
      type_cast_807_inst_ack_1<= rack(0);
      type_cast_807_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_807_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext491_982,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_807_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_824_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_824_inst_req_0;
      type_cast_824_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_824_inst_req_1;
      type_cast_824_inst_ack_1<= rack(0);
      type_cast_824_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_824_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_818,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv156_825,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_840_inst_req_0;
      type_cast_840_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_840_inst_req_1;
      type_cast_840_inst_ack_1<= rack(0);
      type_cast_840_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_840_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call161_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_841,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_861_inst_req_0;
      type_cast_861_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_861_inst_req_1;
      type_cast_861_inst_ack_1<= rack(0);
      type_cast_861_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_861_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_855,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv175_862,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_882_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_882_inst_req_0;
      type_cast_882_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_882_inst_req_1;
      type_cast_882_inst_ack_1<= rack(0);
      type_cast_882_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_882_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call181_876,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_883,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_903_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_903_inst_req_0;
      type_cast_903_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_903_inst_req_1;
      type_cast_903_inst_ack_1<= rack(0);
      type_cast_903_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_903_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call191_897,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv195_904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_924_inst_req_0;
      type_cast_924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_924_inst_req_1;
      type_cast_924_inst_ack_1<= rack(0);
      type_cast_924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call201_918,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_945_inst_req_0;
      type_cast_945_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_945_inst_req_1;
      type_cast_945_inst_ack_1<= rack(0);
      type_cast_945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call211_939,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv215_946,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_966_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_966_inst_req_0;
      type_cast_966_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_966_inst_req_1;
      type_cast_966_inst_ack_1<= rack(0);
      type_cast_966_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_966_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv225_967,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1156_index_1_rename
    process(R_ix_x0x_xlcssa_1155_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1155_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1155_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1156_index_1_resize
    process(ix_x0x_xlcssa_1019) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_1019;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1155_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1156_root_address_inst
    process(array_obj_ref_1156_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1156_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1156_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1309_index_1_rename
    process(R_indvar476_1308_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar476_1308_resized;
      ov(13 downto 0) := iv;
      R_indvar476_1308_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1309_index_1_resize
    process(indvar476_1297) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar476_1297;
      ov := iv(13 downto 0);
      R_indvar476_1308_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1309_root_address_inst
    process(array_obj_ref_1309_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1309_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1309_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1656_index_1_rename
    process(R_ix_x1x_xlcssa_1655_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1655_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1655_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1656_index_1_resize
    process(ix_x1x_xlcssa_1515) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1515;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1655_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1656_root_address_inst
    process(array_obj_ref_1656_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1656_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1656_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_813_index_1_rename
    process(R_indvar490_812_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar490_812_resized;
      ov(13 downto 0) := iv;
      R_indvar490_812_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_813_index_1_resize
    process(indvar490_801) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar490_801;
      ov := iv(13 downto 0);
      R_indvar490_812_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_813_root_address_inst
    process(array_obj_ref_813_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_813_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_813_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_addr_0
    process(ptr_deref_1160_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1160_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1160_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_base_resize
    process(arrayidx237_1158) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx237_1158;
      ov := iv(13 downto 0);
      ptr_deref_1160_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_gather_scatter
    process(shl17x_xi_1151) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl17x_xi_1151;
      ov(63 downto 0) := iv;
      ptr_deref_1160_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_root_address_inst
    process(ptr_deref_1160_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1160_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1160_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1470_addr_0
    process(ptr_deref_1470_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1470_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1470_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1470_base_resize
    process(arrayidx337_1311) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx337_1311;
      ov := iv(13 downto 0);
      ptr_deref_1470_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1470_gather_scatter
    process(add333_1468) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add333_1468;
      ov(63 downto 0) := iv;
      ptr_deref_1470_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1470_root_address_inst
    process(ptr_deref_1470_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1470_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1470_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1660_addr_0
    process(ptr_deref_1660_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1660_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1660_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1660_base_resize
    process(arrayidx352_1658) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx352_1658;
      ov := iv(13 downto 0);
      ptr_deref_1660_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1660_gather_scatter
    process(shl17x_xi436_1651) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl17x_xi436_1651;
      ov(63 downto 0) := iv;
      ptr_deref_1660_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1660_root_address_inst
    process(ptr_deref_1660_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1660_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1660_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_974_addr_0
    process(ptr_deref_974_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_974_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_974_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_974_base_resize
    process(arrayidx_815) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_815;
      ov := iv(13 downto 0);
      ptr_deref_974_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_974_gather_scatter
    process(add226_972) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add226_972;
      ov(63 downto 0) := iv;
      ptr_deref_974_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_974_root_address_inst
    process(ptr_deref_974_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_974_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_974_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1039_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1038;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1039_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1039_branch_req_0,
          ack0 => if_stmt_1039_branch_ack_0,
          ack1 => if_stmt_1039_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1117_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1116;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1117_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1117_branch_req_0,
          ack0 => if_stmt_1117_branch_ack_0,
          ack1 => if_stmt_1117_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1217_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp255443_1216;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1217_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1217_branch_req_0,
          ack0 => if_stmt_1217_branch_ack_0,
          ack1 => if_stmt_1217_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1484_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1483;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1484_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1484_branch_req_0,
          ack0 => if_stmt_1484_branch_ack_0,
          ack1 => if_stmt_1484_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1535_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool344_1534;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1535_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1535_branch_req_0,
          ack0 => if_stmt_1535_branch_ack_0,
          ack1 => if_stmt_1535_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1617_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi428_1616;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1617_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1617_branch_req_0,
          ack0 => if_stmt_1617_branch_ack_0,
          ack1 => if_stmt_1617_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1785_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1784;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1785_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1785_branch_req_0,
          ack0 => if_stmt_1785_branch_ack_0,
          ack1 => if_stmt_1785_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_723_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp447_722;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_723_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_723_branch_req_0,
          ack0 => if_stmt_723_branch_ack_0,
          ack1 => if_stmt_723_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_988_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond32_987;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_988_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_988_branch_req_0,
          ack0 => if_stmt_988_branch_ack_0,
          ack1 => if_stmt_988_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1079_inst
    process(nx_x025x_xi_1060) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x025x_xi_1060, type_cast_1078_wire_constant, tmp_var);
      tmp_1080 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1085_inst
    process(nx_x025x_xi_1060) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x025x_xi_1060, type_cast_1084_wire_constant, tmp_var);
      iNsTr_86_1086 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1579_inst
    process(nx_x025x_xi421_1560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x025x_xi421_1560, type_cast_1578_wire_constant, tmp_var);
      tmp452_1580 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1585_inst
    process(nx_x025x_xi421_1560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x025x_xi421_1560, type_cast_1584_wire_constant, tmp_var);
      iNsTr_134_1586 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1694_inst
    process(add81_599) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add81_599, type_cast_1693_wire_constant, tmp_var);
      sub_1695 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1700_inst
    process(add117_661) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add117_661, type_cast_1699_wire_constant, tmp_var);
      sub395_1701 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1706_inst
    process(add99_630) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add99_630, type_cast_1705_wire_constant, tmp_var);
      tmp453_1707 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1716_inst
    process(tmp3_1711) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1711, type_cast_1715_wire_constant, tmp_var);
      tmp4_1717 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1754_inst
    process(tmp9_1735, mul380_1750) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_1735, mul380_1750, tmp_var);
      mul386_1755 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1778_inst
    process(indvar_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1738, type_cast_1777_wire_constant, tmp_var);
      indvarx_xnext_1779 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1477_inst
    process(indvar476_1297) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar476_1297, type_cast_1476_wire_constant, tmp_var);
      indvarx_xnext477_1478 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_981_inst
    process(indvar490_801) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar490_801, type_cast_980_wire_constant, tmp_var);
      indvarx_xnext491_982 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1056_inst
    process(conv2x_xi_1051) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_1051, type_cast_1055_wire_constant, tmp_var);
      shlx_xi_1057 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1556_inst
    process(conv2x_xi418_1551) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi418_1551, type_cast_1555_wire_constant, tmp_var);
      shlx_xi419_1557 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1031_inst
    process(conv145_716) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv145_716, type_cast_1030_wire_constant, tmp_var);
      and_1032 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1139_inst
    process(Bx_xnot_1134) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1134, type_cast_1138_wire_constant, tmp_var);
      add1519x_xi_1140 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1527_inst
    process(conv249_1210) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv249_1210, type_cast_1526_wire_constant, tmp_var);
      and343_1528 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1639_inst
    process(iNsTr_144_1634) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_144_1634, type_cast_1638_wire_constant, tmp_var);
      add1519x_xi434_1640 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1014_inst
    process(type_cast_1010_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1010_wire, type_cast_1013_wire_constant, tmp_var);
      ASHR_i64_i64_1014_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1208_inst
    process(type_cast_1204_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1204_wire, type_cast_1207_wire_constant, tmp_var);
      ASHR_i64_i64_1208_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1510_inst
    process(type_cast_1506_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1506_wire, type_cast_1509_wire_constant, tmp_var);
      ASHR_i64_i64_1510_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1783_inst
    process(indvarx_xnext_1779, tmp4_1717) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1779, tmp4_1717, tmp_var);
      exitcond5_1784 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1037_inst
    process(and_1032) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_1032, type_cast_1036_wire_constant, tmp_var);
      tobool_1038 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1482_inst
    process(indvarx_xnext477_1478, umax23_1294) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext477_1478, umax23_1294, tmp_var);
      exitcond_1483 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1533_inst
    process(and343_1528) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and343_1528, type_cast_1532_wire_constant, tmp_var);
      tobool344_1534 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_986_inst
    process(indvarx_xnext491_982, umax31_798) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext491_982, umax31_798, tmp_var);
      exitcond32_987 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1228_inst
    process(conv249_1210) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv249_1210, type_cast_1227_wire_constant, tmp_var);
      tmp471_1229 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1280_inst
    process(tmp20_1275) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_1275, type_cast_1279_wire_constant, tmp_var);
      tmp21_1281 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_749_inst
    process(tmp483_744) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp483_744, type_cast_748_wire_constant, tmp_var);
      tmp484_750 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_784_inst
    process(tmp28_779) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp28_779, type_cast_783_wire_constant, tmp_var);
      tmp29_785 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1672_inst
    process(add135_692, add45_537) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add135_692, add45_537, tmp_var);
      mul362_1673 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1677_inst
    process(add81_599, add63_568) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add81_599, add63_568, tmp_var);
      mul375_1678 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1725_inst
    process(add135_692, add45_537) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add135_692, add45_537, tmp_var);
      tmp7_1726 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1734_inst
    process(tmp6_1721, tmp8_1730) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp6_1721, tmp8_1730, tmp_var);
      tmp9_1735 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1749_inst
    process(tmp9_1735, indvar_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_1735, indvar_1738, tmp_var);
      mul380_1750 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_704_inst
    process(conv141_696, add_475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv141_696, add_475, tmp_var);
      mul_705 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_709_inst
    process(mul_705, conv143_700) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_705, conv143_700, tmp_var);
      mul144_710 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_733_inst
    process(add_475, conv141_696) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_475, conv141_696, tmp_var);
      tmp480_734 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_738_inst
    process(tmp480_734, conv143_700) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp480_734, conv143_700, tmp_var);
      tmp482_739 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_764_inst
    process(add_475, tmp24_760) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_475, tmp24_760, tmp_var);
      tmp25_765 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_773_inst
    process(tmp25_765, tmp26_769) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp25_765, tmp26_769, tmp_var);
      tmp27_774 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1184_inst
    process(conv247_1180, conv239_1168) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv247_1180, conv239_1168, tmp_var);
      mul242_1185 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1189_inst
    process(mul242_1185, conv244_1176) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul242_1185, conv244_1176, tmp_var);
      mul245_1190 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1194_inst
    process(mul245_1190, conv241_1172) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul245_1190, conv241_1172, tmp_var);
      mul248_1195 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1247_inst
    process(tmp12_1239, tmp13_1243) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_1239, tmp13_1243, tmp_var);
      tmp14_1248 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1256_inst
    process(tmp14_1248, tmp15_1252) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_1248, tmp15_1252, tmp_var);
      tmp16_1257 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1265_inst
    process(tmp16_1257, tmp17_1261) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_1257, tmp17_1261, tmp_var);
      tmp18_1266 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_505_inst
    process(conv26_501, shl20_491) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv26_501, shl20_491, tmp_var);
      add27_506 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_536_inst
    process(conv44_532, shl38_522) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv44_532, shl38_522, tmp_var);
      add45_537 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_567_inst
    process(conv62_563, shl56_553) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv62_563, shl56_553, tmp_var);
      add63_568 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_598_inst
    process(conv80_594, shl74_584) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv80_594, shl74_584, tmp_var);
      add81_599 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_629_inst
    process(conv98_625, shl92_615) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv98_625, shl92_615, tmp_var);
      add99_630 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_660_inst
    process(conv116_656, shl110_646) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv116_656, shl110_646, tmp_var);
      add117_661 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_691_inst
    process(conv134_687, shl128_677) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv134_687, shl128_677, tmp_var);
      add135_692 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_474_inst
    process(conv9_470, shl_460) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv9_470, shl_460, tmp_var);
      add_475 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1100_inst
    process(conv8x_xi_1096, elementx_x024x_xi_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv8x_xi_1096, elementx_x024x_xi_1067, tmp_var);
      addx_xi_1101 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1341_inst
    process(conv272_1337, shl265_1327) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv272_1337, shl265_1327, tmp_var);
      add273_1342 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1362_inst
    process(shl275_1348, conv282_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl275_1348, conv282_1358, tmp_var);
      add283_1363 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1383_inst
    process(shl285_1369, conv292_1379) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl285_1369, conv292_1379, tmp_var);
      add293_1384 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1404_inst
    process(shl295_1390, conv302_1400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl295_1390, conv302_1400, tmp_var);
      add303_1405 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1425_inst
    process(shl305_1411, conv312_1421) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl305_1411, conv312_1421, tmp_var);
      add313_1426 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1446_inst
    process(shl315_1432, conv322_1442) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl315_1432, conv322_1442, tmp_var);
      add323_1447 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1467_inst
    process(shl325_1453, conv332_1463) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl325_1453, conv332_1463, tmp_var);
      add333_1468 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1600_inst
    process(conv8x_xi424_1596, elementx_x024x_xi422_1567) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv8x_xi424_1596, elementx_x024x_xi422_1567, tmp_var);
      addx_xi425_1601 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_845_inst
    process(conv165_841, shl158_831) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv165_841, shl158_831, tmp_var);
      add166_846 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_866_inst
    process(shl168_852, conv175_862) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_852, conv175_862, tmp_var);
      add176_867 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_887_inst
    process(shl178_873, conv185_883) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl178_873, conv185_883, tmp_var);
      add186_888 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_908_inst
    process(shl188_894, conv195_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl188_894, conv195_904, tmp_var);
      add196_909 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_929_inst
    process(shl198_915, conv205_925) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl198_915, conv205_925, tmp_var);
      add206_930 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_950_inst
    process(shl208_936, conv215_946) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_936, conv215_946, tmp_var);
      add216_951 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_971_inst
    process(shl218_957, conv225_967) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl218_957, conv225_967, tmp_var);
      add226_972 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_490_inst
    process(conv19_485) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_485, type_cast_489_wire_constant, tmp_var);
      shl20_491 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_521_inst
    process(conv37_516) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv37_516, type_cast_520_wire_constant, tmp_var);
      shl38_522 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_552_inst
    process(conv55_547) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv55_547, type_cast_551_wire_constant, tmp_var);
      shl56_553 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_583_inst
    process(conv73_578) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv73_578, type_cast_582_wire_constant, tmp_var);
      shl74_584 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_614_inst
    process(conv91_609) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_609, type_cast_613_wire_constant, tmp_var);
      shl92_615 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_645_inst
    process(conv109_640) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv109_640, type_cast_644_wire_constant, tmp_var);
      shl110_646 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_676_inst
    process(conv127_671) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv127_671, type_cast_675_wire_constant, tmp_var);
      shl128_677 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1050_inst
    process(mul144_710) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul144_710, type_cast_1049_wire_constant, tmp_var);
      conv2x_xi_1051 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_459_inst
    process(conv3_454) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv3_454, type_cast_458_wire_constant, tmp_var);
      shl_460 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1006_inst
    process(umax486_1001) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax486_1001, type_cast_1005_wire_constant, tmp_var);
      tmp487_1007 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1106_inst
    process(addx_xi_1101) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1101, type_cast_1105_wire_constant, tmp_var);
      shl11x_xi_1107 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1133_inst
    process(conv145_716) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv145_716, type_cast_1132_wire_constant, tmp_var);
      Bx_xnot_1134 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1150_inst
    process(shl11x_xix_xlcssa_1124, sh_promx_xi_1146) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl11x_xix_xlcssa_1124, sh_promx_xi_1146, tmp_var);
      shl17x_xi_1151 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1200_inst
    process(mul248_1195) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul248_1195, type_cast_1199_wire_constant, tmp_var);
      sext_1201 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1326_inst
    process(conv263_1321) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv263_1321, type_cast_1325_wire_constant, tmp_var);
      shl265_1327 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1347_inst
    process(add273_1342) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add273_1342, type_cast_1346_wire_constant, tmp_var);
      shl275_1348 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1368_inst
    process(add283_1363) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add283_1363, type_cast_1367_wire_constant, tmp_var);
      shl285_1369 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1389_inst
    process(add293_1384) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add293_1384, type_cast_1388_wire_constant, tmp_var);
      shl295_1390 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1410_inst
    process(add303_1405) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add303_1405, type_cast_1409_wire_constant, tmp_var);
      shl305_1411 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1431_inst
    process(add313_1426) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add313_1426, type_cast_1430_wire_constant, tmp_var);
      shl315_1432 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1452_inst
    process(add323_1447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add323_1447, type_cast_1451_wire_constant, tmp_var);
      shl325_1453 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1502_inst
    process(umax_1497) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1497, type_cast_1501_wire_constant, tmp_var);
      tmp473_1503 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1546_inst
    process(mul248_1195) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul248_1195, type_cast_1545_wire_constant, tmp_var);
      iNsTr_126_1547 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1606_inst
    process(addx_xi425_1601) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi425_1601, type_cast_1605_wire_constant, tmp_var);
      shl11x_xi426_1607 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1633_inst
    process(mul248_1195) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul248_1195, type_cast_1632_wire_constant, tmp_var);
      iNsTr_144_1634 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1650_inst
    process(shl11x_xi426x_xlcssa_1624, sh_promx_xi435_1646) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl11x_xi426x_xlcssa_1624, sh_promx_xi435_1646, tmp_var);
      shl17x_xi436_1651 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_830_inst
    process(conv156_825) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv156_825, type_cast_829_wire_constant, tmp_var);
      shl158_831 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_851_inst
    process(add166_846) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_846, type_cast_850_wire_constant, tmp_var);
      shl168_852 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_872_inst
    process(add176_867) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add176_867, type_cast_871_wire_constant, tmp_var);
      shl178_873 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_893_inst
    process(add186_888) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add186_888, type_cast_892_wire_constant, tmp_var);
      shl188_894 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_914_inst
    process(add196_909) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add196_909, type_cast_913_wire_constant, tmp_var);
      shl198_915 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_935_inst
    process(add206_930) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_930, type_cast_934_wire_constant, tmp_var);
      shl208_936 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_956_inst
    process(add216_951) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add216_951, type_cast_955_wire_constant, tmp_var);
      shl218_957 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1808_inst
    process(conv411_1804, conv356_1796) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv411_1804, conv356_1796, tmp_var);
      sub415_1809 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_721_inst
    process(mul144_710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul144_710, type_cast_720_wire_constant, tmp_var);
      cmp447_722 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1215_inst
    process(conv249_1210) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv249_1210, type_cast_1214_wire_constant, tmp_var);
      cmp255443_1216 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1234_inst
    process(tmp471_1229) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp471_1229, type_cast_1233_wire_constant, tmp_var);
      tmp472_1235 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1286_inst
    process(tmp21_1281) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp21_1281, type_cast_1285_wire_constant, tmp_var);
      tmp22_1287 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_755_inst
    process(tmp484_750) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp484_750, type_cast_754_wire_constant, tmp_var);
      tmp485_756 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_790_inst
    process(tmp29_785) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp29_785, type_cast_789_wire_constant, tmp_var);
      tmp30_791 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1115_inst
    process(convx_xi_1111, shlx_xi_1057) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1111, shlx_xi_1057, tmp_var);
      cmpx_xi_1116 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1615_inst
    process(convx_xi427_1611, shlx_xi419_1557) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi427_1611, shlx_xi419_1557, tmp_var);
      cmpx_xi428_1616 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1145_inst
    process(add1519x_xi_1140) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1519x_xi_1140, type_cast_1144_wire_constant, tmp_var);
      sh_promx_xi_1146 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1645_inst
    process(add1519x_xi434_1640) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1519x_xi434_1640, type_cast_1644_wire_constant, tmp_var);
      sh_promx_xi435_1646 <= tmp_var; --
    end process;
    -- shared split operator group (115) : array_obj_ref_1156_index_offset 
    ApIntAdd_group_115: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1155_scaled;
      array_obj_ref_1156_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1156_index_offset_req_0;
      array_obj_ref_1156_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1156_index_offset_req_1;
      array_obj_ref_1156_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_115_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_115_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_115",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 115
    -- shared split operator group (116) : array_obj_ref_1309_index_offset 
    ApIntAdd_group_116: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar476_1308_scaled;
      array_obj_ref_1309_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1309_index_offset_req_0;
      array_obj_ref_1309_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1309_index_offset_req_1;
      array_obj_ref_1309_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_116_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_116_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_116",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 116
    -- shared split operator group (117) : array_obj_ref_1656_index_offset 
    ApIntAdd_group_117: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1655_scaled;
      array_obj_ref_1656_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1656_index_offset_req_0;
      array_obj_ref_1656_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1656_index_offset_req_1;
      array_obj_ref_1656_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_117_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : array_obj_ref_813_index_offset 
    ApIntAdd_group_118: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar490_812_scaled;
      array_obj_ref_813_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_813_index_offset_req_0;
      array_obj_ref_813_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_813_index_offset_req_1;
      array_obj_ref_813_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_118_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- unary operator type_cast_1273_inst
    process(tmp19_1270) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp19_1270, tmp_var);
      type_cast_1273_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1794_inst
    process(call355_1667) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call355_1667, tmp_var);
      type_cast_1794_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1802_inst
    process(call410_1799) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call410_1799, tmp_var);
      type_cast_1802_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_714_inst
    process(mul144_710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul144_710, tmp_var);
      type_cast_714_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_742_inst
    process(tmp482_739) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp482_739, tmp_var);
      type_cast_742_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_777_inst
    process(tmp27_774) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp27_774, tmp_var);
      type_cast_777_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_974_store_0 ptr_deref_1160_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_974_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1160_store_0_req_0;
      ptr_deref_974_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1160_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_974_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1160_store_0_req_1;
      ptr_deref_974_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1160_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_974_word_address_0 & ptr_deref_1160_word_address_0;
      data_in <= ptr_deref_974_data_0 & ptr_deref_1160_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1470_store_0 ptr_deref_1660_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1470_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1660_store_0_req_0;
      ptr_deref_1470_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1660_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1470_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1660_store_0_req_1;
      ptr_deref_1470_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1660_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1470_word_address_0 & ptr_deref_1660_word_address_0;
      data_in <= ptr_deref_1470_data_0 & ptr_deref_1660_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_938_inst RPIPE_maxpool_input_pipe_1313_inst RPIPE_maxpool_input_pipe_875_inst RPIPE_maxpool_input_pipe_1392_inst RPIPE_maxpool_input_pipe_817_inst RPIPE_maxpool_input_pipe_1329_inst RPIPE_maxpool_input_pipe_959_inst RPIPE_maxpool_input_pipe_1455_inst RPIPE_maxpool_input_pipe_896_inst RPIPE_maxpool_input_pipe_1088_inst RPIPE_maxpool_input_pipe_1350_inst RPIPE_maxpool_input_pipe_833_inst RPIPE_maxpool_input_pipe_1413_inst RPIPE_maxpool_input_pipe_854_inst RPIPE_maxpool_input_pipe_1434_inst RPIPE_maxpool_input_pipe_917_inst RPIPE_maxpool_input_pipe_1371_inst RPIPE_maxpool_input_pipe_446_inst RPIPE_maxpool_input_pipe_462_inst RPIPE_maxpool_input_pipe_477_inst RPIPE_maxpool_input_pipe_493_inst RPIPE_maxpool_input_pipe_508_inst RPIPE_maxpool_input_pipe_524_inst RPIPE_maxpool_input_pipe_539_inst RPIPE_maxpool_input_pipe_555_inst RPIPE_maxpool_input_pipe_570_inst RPIPE_maxpool_input_pipe_586_inst RPIPE_maxpool_input_pipe_601_inst RPIPE_maxpool_input_pipe_617_inst RPIPE_maxpool_input_pipe_632_inst RPIPE_maxpool_input_pipe_648_inst RPIPE_maxpool_input_pipe_663_inst RPIPE_maxpool_input_pipe_679_inst RPIPE_maxpool_input_pipe_1588_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_938_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_1313_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_875_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_1392_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_817_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_1329_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_959_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_1455_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_896_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_1088_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_1350_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_833_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_1413_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_854_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_1434_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_917_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_1371_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_446_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_462_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_477_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_493_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_508_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_524_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_539_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_555_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_570_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_586_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_601_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_617_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_632_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_648_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_663_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_679_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1588_inst_req_0;
      RPIPE_maxpool_input_pipe_938_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_1313_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_875_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_1392_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_817_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_1329_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_959_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_1455_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_896_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_1088_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_1350_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_833_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_1413_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_854_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_1434_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_917_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_1371_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_446_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_462_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_477_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_493_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_508_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_524_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_539_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_555_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_570_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_586_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_601_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_617_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_632_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_648_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_663_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_679_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1588_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_938_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_1313_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_875_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_1392_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_817_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_1329_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_959_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_1455_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_896_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_1088_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_1350_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_833_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_1413_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_854_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_1434_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_917_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_1371_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_446_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_462_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_477_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_493_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_508_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_524_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_539_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_555_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_570_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_586_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_601_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_617_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_632_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_648_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_663_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_679_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1588_inst_req_1;
      RPIPE_maxpool_input_pipe_938_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_1313_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_875_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_1392_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_817_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_1329_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_959_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_1455_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_896_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_1088_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_1350_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_833_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_1413_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_854_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_1434_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_917_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_1371_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_446_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_462_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_477_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_493_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_508_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_524_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_539_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_555_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_570_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_586_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_601_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_617_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_632_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_648_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_663_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_679_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1588_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call211_939 <= data_out(271 downto 264);
      call260_1314 <= data_out(263 downto 256);
      call181_876 <= data_out(255 downto 248);
      call298_1393 <= data_out(247 downto 240);
      call153_818 <= data_out(239 downto 232);
      call268_1330 <= data_out(231 downto 224);
      call221_960 <= data_out(223 downto 216);
      call328_1456 <= data_out(215 downto 208);
      call191_897 <= data_out(207 downto 200);
      callx_xi_1089 <= data_out(199 downto 192);
      call278_1351 <= data_out(191 downto 184);
      call161_834 <= data_out(183 downto 176);
      call308_1414 <= data_out(175 downto 168);
      call171_855 <= data_out(167 downto 160);
      call318_1435 <= data_out(159 downto 152);
      call201_918 <= data_out(151 downto 144);
      call288_1372 <= data_out(143 downto 136);
      call_447 <= data_out(135 downto 128);
      call6_463 <= data_out(127 downto 120);
      call14_478 <= data_out(119 downto 112);
      call23_494 <= data_out(111 downto 104);
      call32_509 <= data_out(103 downto 96);
      call41_525 <= data_out(95 downto 88);
      call50_540 <= data_out(87 downto 80);
      call59_556 <= data_out(79 downto 72);
      call68_571 <= data_out(71 downto 64);
      call77_587 <= data_out(63 downto 56);
      call86_602 <= data_out(55 downto 48);
      call95_618 <= data_out(47 downto 40);
      call104_633 <= data_out(39 downto 32);
      call113_649 <= data_out(31 downto 24);
      call122_664 <= data_out(23 downto 16);
      call131_680 <= data_out(15 downto 8);
      callx_xi423_1589 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1810_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1810_inst_req_0;
      WPIPE_elapsed_time_pipe_1810_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1810_inst_req_1;
      WPIPE_elapsed_time_pipe_1810_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub415_1809;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_maxpool_output_pipe_1090_inst WPIPE_maxpool_output_pipe_940_inst WPIPE_maxpool_output_pipe_1373_inst WPIPE_maxpool_output_pipe_919_inst WPIPE_maxpool_output_pipe_1315_inst WPIPE_maxpool_output_pipe_1394_inst WPIPE_maxpool_output_pipe_819_inst WPIPE_maxpool_output_pipe_1331_inst WPIPE_maxpool_output_pipe_961_inst WPIPE_maxpool_output_pipe_1436_inst WPIPE_maxpool_output_pipe_1415_inst WPIPE_maxpool_output_pipe_877_inst WPIPE_maxpool_output_pipe_835_inst WPIPE_maxpool_output_pipe_1352_inst WPIPE_maxpool_output_pipe_856_inst WPIPE_maxpool_output_pipe_1457_inst WPIPE_maxpool_output_pipe_898_inst WPIPE_maxpool_output_pipe_437_inst WPIPE_maxpool_output_pipe_441_inst WPIPE_maxpool_output_pipe_448_inst WPIPE_maxpool_output_pipe_464_inst WPIPE_maxpool_output_pipe_479_inst WPIPE_maxpool_output_pipe_495_inst WPIPE_maxpool_output_pipe_510_inst WPIPE_maxpool_output_pipe_526_inst WPIPE_maxpool_output_pipe_541_inst WPIPE_maxpool_output_pipe_557_inst WPIPE_maxpool_output_pipe_572_inst WPIPE_maxpool_output_pipe_588_inst WPIPE_maxpool_output_pipe_603_inst WPIPE_maxpool_output_pipe_619_inst WPIPE_maxpool_output_pipe_634_inst WPIPE_maxpool_output_pipe_650_inst WPIPE_maxpool_output_pipe_665_inst WPIPE_maxpool_output_pipe_681_inst WPIPE_maxpool_output_pipe_1590_inst WPIPE_maxpool_output_pipe_1682_inst WPIPE_maxpool_output_pipe_1686_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(303 downto 0);
      signal sample_req, sample_ack : BooleanArray( 37 downto 0);
      signal update_req, update_ack : BooleanArray( 37 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 37 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 37 downto 0);
      signal guard_vector : std_logic_vector( 37 downto 0);
      constant inBUFs : IntegerArray(37 downto 0) := (37 => 0, 36 => 0, 35 => 0, 34 => 0, 33 => 0, 32 => 0, 31 => 0, 30 => 0, 29 => 0, 28 => 0, 27 => 0, 26 => 0, 25 => 0, 24 => 0, 23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(37 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false);
      constant guardBuffering: IntegerArray(37 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2);
      -- 
    begin -- 
      sample_req_unguarded(37) <= WPIPE_maxpool_output_pipe_1090_inst_req_0;
      sample_req_unguarded(36) <= WPIPE_maxpool_output_pipe_940_inst_req_0;
      sample_req_unguarded(35) <= WPIPE_maxpool_output_pipe_1373_inst_req_0;
      sample_req_unguarded(34) <= WPIPE_maxpool_output_pipe_919_inst_req_0;
      sample_req_unguarded(33) <= WPIPE_maxpool_output_pipe_1315_inst_req_0;
      sample_req_unguarded(32) <= WPIPE_maxpool_output_pipe_1394_inst_req_0;
      sample_req_unguarded(31) <= WPIPE_maxpool_output_pipe_819_inst_req_0;
      sample_req_unguarded(30) <= WPIPE_maxpool_output_pipe_1331_inst_req_0;
      sample_req_unguarded(29) <= WPIPE_maxpool_output_pipe_961_inst_req_0;
      sample_req_unguarded(28) <= WPIPE_maxpool_output_pipe_1436_inst_req_0;
      sample_req_unguarded(27) <= WPIPE_maxpool_output_pipe_1415_inst_req_0;
      sample_req_unguarded(26) <= WPIPE_maxpool_output_pipe_877_inst_req_0;
      sample_req_unguarded(25) <= WPIPE_maxpool_output_pipe_835_inst_req_0;
      sample_req_unguarded(24) <= WPIPE_maxpool_output_pipe_1352_inst_req_0;
      sample_req_unguarded(23) <= WPIPE_maxpool_output_pipe_856_inst_req_0;
      sample_req_unguarded(22) <= WPIPE_maxpool_output_pipe_1457_inst_req_0;
      sample_req_unguarded(21) <= WPIPE_maxpool_output_pipe_898_inst_req_0;
      sample_req_unguarded(20) <= WPIPE_maxpool_output_pipe_437_inst_req_0;
      sample_req_unguarded(19) <= WPIPE_maxpool_output_pipe_441_inst_req_0;
      sample_req_unguarded(18) <= WPIPE_maxpool_output_pipe_448_inst_req_0;
      sample_req_unguarded(17) <= WPIPE_maxpool_output_pipe_464_inst_req_0;
      sample_req_unguarded(16) <= WPIPE_maxpool_output_pipe_479_inst_req_0;
      sample_req_unguarded(15) <= WPIPE_maxpool_output_pipe_495_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_maxpool_output_pipe_510_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_maxpool_output_pipe_526_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_maxpool_output_pipe_541_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_maxpool_output_pipe_557_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_maxpool_output_pipe_572_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_588_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_603_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_619_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_634_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_650_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_665_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_681_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1590_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1682_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1686_inst_req_0;
      WPIPE_maxpool_output_pipe_1090_inst_ack_0 <= sample_ack_unguarded(37);
      WPIPE_maxpool_output_pipe_940_inst_ack_0 <= sample_ack_unguarded(36);
      WPIPE_maxpool_output_pipe_1373_inst_ack_0 <= sample_ack_unguarded(35);
      WPIPE_maxpool_output_pipe_919_inst_ack_0 <= sample_ack_unguarded(34);
      WPIPE_maxpool_output_pipe_1315_inst_ack_0 <= sample_ack_unguarded(33);
      WPIPE_maxpool_output_pipe_1394_inst_ack_0 <= sample_ack_unguarded(32);
      WPIPE_maxpool_output_pipe_819_inst_ack_0 <= sample_ack_unguarded(31);
      WPIPE_maxpool_output_pipe_1331_inst_ack_0 <= sample_ack_unguarded(30);
      WPIPE_maxpool_output_pipe_961_inst_ack_0 <= sample_ack_unguarded(29);
      WPIPE_maxpool_output_pipe_1436_inst_ack_0 <= sample_ack_unguarded(28);
      WPIPE_maxpool_output_pipe_1415_inst_ack_0 <= sample_ack_unguarded(27);
      WPIPE_maxpool_output_pipe_877_inst_ack_0 <= sample_ack_unguarded(26);
      WPIPE_maxpool_output_pipe_835_inst_ack_0 <= sample_ack_unguarded(25);
      WPIPE_maxpool_output_pipe_1352_inst_ack_0 <= sample_ack_unguarded(24);
      WPIPE_maxpool_output_pipe_856_inst_ack_0 <= sample_ack_unguarded(23);
      WPIPE_maxpool_output_pipe_1457_inst_ack_0 <= sample_ack_unguarded(22);
      WPIPE_maxpool_output_pipe_898_inst_ack_0 <= sample_ack_unguarded(21);
      WPIPE_maxpool_output_pipe_437_inst_ack_0 <= sample_ack_unguarded(20);
      WPIPE_maxpool_output_pipe_441_inst_ack_0 <= sample_ack_unguarded(19);
      WPIPE_maxpool_output_pipe_448_inst_ack_0 <= sample_ack_unguarded(18);
      WPIPE_maxpool_output_pipe_464_inst_ack_0 <= sample_ack_unguarded(17);
      WPIPE_maxpool_output_pipe_479_inst_ack_0 <= sample_ack_unguarded(16);
      WPIPE_maxpool_output_pipe_495_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_maxpool_output_pipe_510_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_maxpool_output_pipe_526_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_maxpool_output_pipe_541_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_maxpool_output_pipe_557_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_maxpool_output_pipe_572_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_maxpool_output_pipe_588_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_603_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_619_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_634_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_650_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_665_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_681_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1590_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1682_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1686_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(37) <= WPIPE_maxpool_output_pipe_1090_inst_req_1;
      update_req_unguarded(36) <= WPIPE_maxpool_output_pipe_940_inst_req_1;
      update_req_unguarded(35) <= WPIPE_maxpool_output_pipe_1373_inst_req_1;
      update_req_unguarded(34) <= WPIPE_maxpool_output_pipe_919_inst_req_1;
      update_req_unguarded(33) <= WPIPE_maxpool_output_pipe_1315_inst_req_1;
      update_req_unguarded(32) <= WPIPE_maxpool_output_pipe_1394_inst_req_1;
      update_req_unguarded(31) <= WPIPE_maxpool_output_pipe_819_inst_req_1;
      update_req_unguarded(30) <= WPIPE_maxpool_output_pipe_1331_inst_req_1;
      update_req_unguarded(29) <= WPIPE_maxpool_output_pipe_961_inst_req_1;
      update_req_unguarded(28) <= WPIPE_maxpool_output_pipe_1436_inst_req_1;
      update_req_unguarded(27) <= WPIPE_maxpool_output_pipe_1415_inst_req_1;
      update_req_unguarded(26) <= WPIPE_maxpool_output_pipe_877_inst_req_1;
      update_req_unguarded(25) <= WPIPE_maxpool_output_pipe_835_inst_req_1;
      update_req_unguarded(24) <= WPIPE_maxpool_output_pipe_1352_inst_req_1;
      update_req_unguarded(23) <= WPIPE_maxpool_output_pipe_856_inst_req_1;
      update_req_unguarded(22) <= WPIPE_maxpool_output_pipe_1457_inst_req_1;
      update_req_unguarded(21) <= WPIPE_maxpool_output_pipe_898_inst_req_1;
      update_req_unguarded(20) <= WPIPE_maxpool_output_pipe_437_inst_req_1;
      update_req_unguarded(19) <= WPIPE_maxpool_output_pipe_441_inst_req_1;
      update_req_unguarded(18) <= WPIPE_maxpool_output_pipe_448_inst_req_1;
      update_req_unguarded(17) <= WPIPE_maxpool_output_pipe_464_inst_req_1;
      update_req_unguarded(16) <= WPIPE_maxpool_output_pipe_479_inst_req_1;
      update_req_unguarded(15) <= WPIPE_maxpool_output_pipe_495_inst_req_1;
      update_req_unguarded(14) <= WPIPE_maxpool_output_pipe_510_inst_req_1;
      update_req_unguarded(13) <= WPIPE_maxpool_output_pipe_526_inst_req_1;
      update_req_unguarded(12) <= WPIPE_maxpool_output_pipe_541_inst_req_1;
      update_req_unguarded(11) <= WPIPE_maxpool_output_pipe_557_inst_req_1;
      update_req_unguarded(10) <= WPIPE_maxpool_output_pipe_572_inst_req_1;
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_588_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_603_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_619_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_634_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_650_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_665_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_681_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1590_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1682_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1686_inst_req_1;
      WPIPE_maxpool_output_pipe_1090_inst_ack_1 <= update_ack_unguarded(37);
      WPIPE_maxpool_output_pipe_940_inst_ack_1 <= update_ack_unguarded(36);
      WPIPE_maxpool_output_pipe_1373_inst_ack_1 <= update_ack_unguarded(35);
      WPIPE_maxpool_output_pipe_919_inst_ack_1 <= update_ack_unguarded(34);
      WPIPE_maxpool_output_pipe_1315_inst_ack_1 <= update_ack_unguarded(33);
      WPIPE_maxpool_output_pipe_1394_inst_ack_1 <= update_ack_unguarded(32);
      WPIPE_maxpool_output_pipe_819_inst_ack_1 <= update_ack_unguarded(31);
      WPIPE_maxpool_output_pipe_1331_inst_ack_1 <= update_ack_unguarded(30);
      WPIPE_maxpool_output_pipe_961_inst_ack_1 <= update_ack_unguarded(29);
      WPIPE_maxpool_output_pipe_1436_inst_ack_1 <= update_ack_unguarded(28);
      WPIPE_maxpool_output_pipe_1415_inst_ack_1 <= update_ack_unguarded(27);
      WPIPE_maxpool_output_pipe_877_inst_ack_1 <= update_ack_unguarded(26);
      WPIPE_maxpool_output_pipe_835_inst_ack_1 <= update_ack_unguarded(25);
      WPIPE_maxpool_output_pipe_1352_inst_ack_1 <= update_ack_unguarded(24);
      WPIPE_maxpool_output_pipe_856_inst_ack_1 <= update_ack_unguarded(23);
      WPIPE_maxpool_output_pipe_1457_inst_ack_1 <= update_ack_unguarded(22);
      WPIPE_maxpool_output_pipe_898_inst_ack_1 <= update_ack_unguarded(21);
      WPIPE_maxpool_output_pipe_437_inst_ack_1 <= update_ack_unguarded(20);
      WPIPE_maxpool_output_pipe_441_inst_ack_1 <= update_ack_unguarded(19);
      WPIPE_maxpool_output_pipe_448_inst_ack_1 <= update_ack_unguarded(18);
      WPIPE_maxpool_output_pipe_464_inst_ack_1 <= update_ack_unguarded(17);
      WPIPE_maxpool_output_pipe_479_inst_ack_1 <= update_ack_unguarded(16);
      WPIPE_maxpool_output_pipe_495_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_maxpool_output_pipe_510_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_maxpool_output_pipe_526_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_maxpool_output_pipe_541_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_maxpool_output_pipe_557_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_maxpool_output_pipe_572_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_maxpool_output_pipe_588_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_603_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_619_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_634_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_650_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_665_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_681_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1590_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1682_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1686_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      data_in <= callx_xi_1089 & call211_939 & call288_1372 & call201_918 & call260_1314 & call298_1393 & call153_818 & call268_1330 & call221_960 & call318_1435 & call308_1414 & call181_876 & call161_834 & call278_1351 & call171_855 & call328_1456 & call191_897 & type_cast_439_wire_constant & type_cast_443_wire_constant & call_447 & call6_463 & call14_478 & call23_494 & call32_509 & call41_525 & call50_540 & call59_556 & call68_571 & call77_587 & call86_602 & call95_618 & call104_633 & call113_649 & call122_664 & call131_680 & callx_xi423_1589 & type_cast_1684_wire_constant & type_cast_1688_wire_constant;
      maxpool_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_1_gI", nreqs => 38, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 38, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_num_out_pipe_1679_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1679_inst_req_0;
      WPIPE_num_out_pipe_1679_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1679_inst_req_1;
      WPIPE_num_out_pipe_1679_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= mul375_1678;
      num_out_pipe_write_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_1667_call call_stmt_1799_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1667_call_req_0;
      reqL_unguarded(0) <= call_stmt_1799_call_req_0;
      call_stmt_1667_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1799_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1667_call_req_1;
      reqR_unguarded(0) <= call_stmt_1799_call_req_1;
      call_stmt_1667_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1799_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call355_1667 <= data_out(127 downto 64);
      call410_1799 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1766_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1766_call_req_0;
      call_stmt_1766_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1766_call_req_1;
      call_stmt_1766_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv381_1759 & conv387_1763;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(127 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1773_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1773_call_req_0;
      call_stmt_1773_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1773_call_req_1;
      call_stmt_1773_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul362_1673 & add63_568 & sub_1695 & sub395_1701 & add45_537 & add27_506;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(95 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_4332_start: Boolean;
  signal convolve_CP_4332_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1845_req_0 : boolean;
  signal RPIPE_kernel_pipe1_1859_inst_req_0 : boolean;
  signal phi_stmt_1845_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1859_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1907_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_1907_inst_ack_1 : boolean;
  signal RPIPE_input_pipe1_1852_inst_ack_0 : boolean;
  signal phi_stmt_1845_req_1 : boolean;
  signal n_out_count_1921_1849_buf_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1907_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_1907_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1943_inst_req_0 : boolean;
  signal n_out_count_1921_1849_buf_req_1 : boolean;
  signal SUB_u32_u32_1873_inst_req_0 : boolean;
  signal SUB_u32_u32_1873_inst_ack_0 : boolean;
  signal slice_1937_inst_req_1 : boolean;
  signal nacc_1892_1843_buf_req_0 : boolean;
  signal W_next_sum_1915_delayed_1_0_1939_inst_req_0 : boolean;
  signal slice_1937_inst_ack_1 : boolean;
  signal type_cast_1945_inst_req_0 : boolean;
  signal nacc_1892_1843_buf_ack_0 : boolean;
  signal n_out_count_1921_1849_buf_ack_1 : boolean;
  signal type_cast_1945_inst_ack_0 : boolean;
  signal SUB_u32_u32_1873_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_1928_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_1928_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1943_inst_ack_0 : boolean;
  signal SUB_u32_u32_1873_inst_ack_1 : boolean;
  signal slice_1937_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_1852_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1943_inst_req_1 : boolean;
  signal W_next_sum_1915_delayed_1_0_1939_inst_req_1 : boolean;
  signal type_cast_1945_inst_ack_1 : boolean;
  signal nacc_1892_1843_buf_req_1 : boolean;
  signal nacc_1892_1843_buf_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_1859_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_1928_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_1852_inst_ack_1 : boolean;
  signal W_next_sum_1915_delayed_1_0_1939_inst_ack_1 : boolean;
  signal n_out_count_1921_1849_buf_req_0 : boolean;
  signal slice_1933_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_1928_inst_ack_1 : boolean;
  signal slice_1933_inst_req_1 : boolean;
  signal slice_1933_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_1852_inst_req_0 : boolean;
  signal W_next_sum_1915_delayed_1_0_1939_inst_ack_0 : boolean;
  signal slice_1933_inst_ack_1 : boolean;
  signal type_cast_1945_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_1859_inst_ack_1 : boolean;
  signal slice_1937_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1821_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1821_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1821_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1821_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1824_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1824_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1824_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1824_inst_ack_1 : boolean;
  signal do_while_stmt_1835_branch_req_0 : boolean;
  signal phi_stmt_1837_req_0 : boolean;
  signal phi_stmt_1837_req_1 : boolean;
  signal phi_stmt_1837_ack_0 : boolean;
  signal nmycount_1900_1839_buf_req_0 : boolean;
  signal nmycount_1900_1839_buf_ack_0 : boolean;
  signal nmycount_1900_1839_buf_req_1 : boolean;
  signal nmycount_1900_1839_buf_ack_1 : boolean;
  signal phi_stmt_1841_req_0 : boolean;
  signal phi_stmt_1841_req_1 : boolean;
  signal phi_stmt_1841_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1943_inst_ack_1 : boolean;
  signal W_next_sum_1920_delayed_1_0_1947_inst_req_0 : boolean;
  signal W_next_sum_1920_delayed_1_0_1947_inst_ack_0 : boolean;
  signal W_next_sum_1920_delayed_1_0_1947_inst_req_1 : boolean;
  signal W_next_sum_1920_delayed_1_0_1947_inst_ack_1 : boolean;
  signal type_cast_1953_inst_req_0 : boolean;
  signal type_cast_1953_inst_ack_0 : boolean;
  signal type_cast_1953_inst_req_1 : boolean;
  signal type_cast_1953_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1951_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1951_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1951_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1951_inst_ack_1 : boolean;
  signal do_while_stmt_1835_branch_ack_0 : boolean;
  signal do_while_stmt_1835_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_4332_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4332_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_4332_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4332_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_4332: Block -- control-path 
    signal convolve_CP_4332_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convolve_CP_4332_elements(0) <= convolve_CP_4332_start;
    convolve_CP_4332_symbol <= convolve_CP_4332_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1819/$entry
      -- CP-element group 0: 	 branch_block_stmt_1819/branch_block_stmt_1819__entry__
      -- CP-element group 0: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834__entry__
      -- CP-element group 0: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/$entry
      -- CP-element group 0: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_Sample/rr
      -- 
    rr_4354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(0), ack => RPIPE_num_out_pipe_1821_inst_req_0); -- 
    rr_4368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(0), ack => RPIPE_size_pipe_1824_inst_req_0); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1819/$exit
      -- CP-element group 1: 	 branch_block_stmt_1819/branch_block_stmt_1819__exit__
      -- CP-element group 1: 	 branch_block_stmt_1819/do_while_stmt_1835__exit__
      -- 
    convolve_CP_4332_elements(1) <= convolve_CP_4332_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_Update/cr
      -- 
    ra_4355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1821_inst_ack_0, ack => convolve_CP_4332_elements(2)); -- 
    cr_4359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(2), ack => RPIPE_num_out_pipe_1821_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_num_out_pipe_1821_Update/ca
      -- 
    ca_4360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1821_inst_ack_1, ack => convolve_CP_4332_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_Update/cr
      -- 
    ra_4369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1824_inst_ack_0, ack => convolve_CP_4332_elements(4)); -- 
    cr_4373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(4), ack => RPIPE_size_pipe_1824_inst_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/RPIPE_size_pipe_1824_Update/ca
      -- 
    ca_4374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1824_inst_ack_1, ack => convolve_CP_4332_elements(5)); -- 
    -- CP-element group 6:  join  transition  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834__exit__
      -- CP-element group 6: 	 branch_block_stmt_1819/do_while_stmt_1835__entry__
      -- CP-element group 6: 	 branch_block_stmt_1819/assign_stmt_1822_to_assign_stmt_1834/$exit
      -- 
    convolve_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "convolve_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(3) & convolve_CP_4332_elements(5);
      gj_convolve_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1819/do_while_stmt_1835/$entry
      -- CP-element group 7: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835__entry__
      -- 
    convolve_CP_4332_elements(7) <= convolve_CP_4332_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	127 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835__exit__
      -- 
    -- Element group convolve_CP_4332_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1819/do_while_stmt_1835/loop_back
      -- 
    -- Element group convolve_CP_4332_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	125 
    -- CP-element group 10: 	126 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1819/do_while_stmt_1835/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1819/do_while_stmt_1835/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1819/do_while_stmt_1835/loop_taken/$entry
      -- 
    convolve_CP_4332_elements(10) <= convolve_CP_4332_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	124 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1819/do_while_stmt_1835/loop_body_done
      -- 
    convolve_CP_4332_elements(11) <= convolve_CP_4332_elements(124);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	62 
    -- CP-element group 12: 	45 
    -- CP-element group 12: 	26 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_4332_elements(12) <= convolve_CP_4332_elements(9);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	64 
    -- CP-element group 13: 	47 
    -- CP-element group 13: 	28 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_4332_elements(13) <= convolve_CP_4332_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	83 
    -- CP-element group 14: 	123 
    -- CP-element group 14: 	58 
    -- CP-element group 14: 	59 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	21 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	40 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_4332_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	123 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/condition_evaluated
      -- 
    condition_evaluated_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(15), ack => do_while_stmt_1835_branch_req_0); -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(123) & convolve_CP_4332_elements(19);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	39 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_sample_start__ps
      -- CP-element group 16: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/aggregated_phi_sample_req
      -- 
    convolve_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(58) & convolve_CP_4332_elements(20) & convolve_CP_4332_elements(39) & convolve_CP_4332_elements(19);
      gj_convolve_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	60 
    -- CP-element group 17: 	42 
    -- CP-element group 17: 	23 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	76 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	84 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	58 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	39 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_sample_completed_
      -- 
    convolve_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(60) & convolve_CP_4332_elements(42) & convolve_CP_4332_elements(23);
      gj_convolve_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	40 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	43 
    -- CP-element group 18: 	24 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_update_start__ps
      -- CP-element group 18: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/aggregated_phi_update_req
      -- 
    convolve_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(59) & convolve_CP_4332_elements(21) & convolve_CP_4332_elements(40);
      gj_convolve_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	61 
    -- CP-element group 19: 	44 
    -- CP-element group 19: 	25 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(61) & convolve_CP_4332_elements(44) & convolve_CP_4332_elements(25);
      gj_convolve_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	86 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_sample_start_
      -- 
    convolve_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(86) & convolve_CP_4332_elements(17);
      gj_convolve_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	91 
    -- CP-element group 21: 	114 
    -- CP-element group 21: 	103 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_update_start_
      -- 
    convolve_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(91) & convolve_CP_4332_elements(114) & convolve_CP_4332_elements(103);
      gj_convolve_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_sample_start__ps
      -- 
    convolve_CP_4332_elements(22) <= convolve_CP_4332_elements(16);
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	17 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_sample_completed__ps
      -- 
    -- Element group convolve_CP_4332_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_update_start__ps
      -- 
    convolve_CP_4332_elements(24) <= convolve_CP_4332_elements(18);
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	90 
    -- CP-element group 25: 	112 
    -- CP-element group 25: 	101 
    -- CP-element group 25: 	19 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_update_completed__ps
      -- 
    -- Element group convolve_CP_4332_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	12 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_loopback_trigger
      -- 
    convolve_CP_4332_elements(26) <= convolve_CP_4332_elements(12);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_loopback_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_loopback_sample_req_ps
      -- 
    phi_stmt_1837_loopback_sample_req_4404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1837_loopback_sample_req_4404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(27), ack => phi_stmt_1837_req_0); -- 
    -- Element group convolve_CP_4332_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	13 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_entry_trigger
      -- 
    convolve_CP_4332_elements(28) <= convolve_CP_4332_elements(13);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_entry_sample_req
      -- CP-element group 29: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_entry_sample_req_ps
      -- 
    phi_stmt_1837_entry_sample_req_4407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1837_entry_sample_req_4407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(29), ack => phi_stmt_1837_req_1); -- 
    -- Element group convolve_CP_4332_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_phi_mux_ack
      -- CP-element group 30: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1837_phi_mux_ack_ps
      -- 
    phi_stmt_1837_phi_mux_ack_4410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1837_ack_0, ack => convolve_CP_4332_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_Sample/req
      -- 
    req_4423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(31), ack => nmycount_1900_1839_buf_req_0); -- 
    -- Element group convolve_CP_4332_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_Update/req
      -- 
    req_4428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(32), ack => nmycount_1900_1839_buf_req_1); -- 
    -- Element group convolve_CP_4332_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_Sample/ack
      -- 
    ack_4424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1900_1839_buf_ack_0, ack => convolve_CP_4332_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_update_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nmycount_1839_Update/ack
      -- 
    ack_4429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1900_1839_buf_ack_1, ack => convolve_CP_4332_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_mcount_var_1840_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_mcount_var_1840_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_mcount_var_1840_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_mcount_var_1840_sample_completed_
      -- 
    -- Element group convolve_CP_4332_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_mcount_var_1840_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_mcount_var_1840_update_start_
      -- 
    -- Element group convolve_CP_4332_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_mcount_var_1840_update_completed__ps
      -- 
    convolve_CP_4332_elements(37) <= convolve_CP_4332_elements(38);
    -- CP-element group 38:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	37 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_mcount_var_1840_update_completed_
      -- 
    -- Element group convolve_CP_4332_elements(38) is a control-delay.
    cp_element_38_delay: control_delay_element  generic map(name => " 38_delay", delay_value => 1)  port map(req => convolve_CP_4332_elements(36), ack => convolve_CP_4332_elements(38), clk => clk, reset =>reset);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	86 
    -- CP-element group 39: 	78 
    -- CP-element group 39: 	82 
    -- CP-element group 39: 	17 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	16 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_sample_start_
      -- 
    convolve_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(86) & convolve_CP_4332_elements(78) & convolve_CP_4332_elements(82) & convolve_CP_4332_elements(17);
      gj_convolve_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	14 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	95 
    -- CP-element group 40: 	99 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	18 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_update_start_
      -- 
    convolve_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(95) & convolve_CP_4332_elements(99);
      gj_convolve_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_sample_start__ps
      -- 
    convolve_CP_4332_elements(41) <= convolve_CP_4332_elements(16);
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	17 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_sample_completed__ps
      -- 
    -- Element group convolve_CP_4332_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	18 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_update_start__ps
      -- 
    convolve_CP_4332_elements(43) <= convolve_CP_4332_elements(18);
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	93 
    -- CP-element group 44: 	97 
    -- CP-element group 44: 	19 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_update_completed__ps
      -- 
    -- Element group convolve_CP_4332_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	12 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_loopback_trigger
      -- 
    convolve_CP_4332_elements(45) <= convolve_CP_4332_elements(12);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_loopback_sample_req
      -- CP-element group 46: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_loopback_sample_req_ps
      -- 
    phi_stmt_1841_loopback_sample_req_4448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1841_loopback_sample_req_4448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(46), ack => phi_stmt_1841_req_0); -- 
    -- Element group convolve_CP_4332_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	13 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_entry_trigger
      -- 
    convolve_CP_4332_elements(47) <= convolve_CP_4332_elements(13);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_entry_sample_req
      -- CP-element group 48: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_entry_sample_req_ps
      -- 
    phi_stmt_1841_entry_sample_req_4451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1841_entry_sample_req_4451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(48), ack => phi_stmt_1841_req_1); -- 
    -- Element group convolve_CP_4332_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_phi_mux_ack
      -- CP-element group 49: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1841_phi_mux_ack_ps
      -- 
    phi_stmt_1841_phi_mux_ack_4454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1841_ack_0, ack => convolve_CP_4332_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_Sample/req
      -- CP-element group 50: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_sample_start__ps
      -- 
    req_4467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(50), ack => nacc_1892_1843_buf_req_0); -- 
    -- Element group convolve_CP_4332_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_Update/req
      -- CP-element group 51: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_update_start__ps
      -- 
    req_4472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(51), ack => nacc_1892_1843_buf_req_1); -- 
    -- Element group convolve_CP_4332_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_sample_completed__ps
      -- 
    ack_4468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1892_1843_buf_ack_0, ack => convolve_CP_4332_elements(52)); -- 
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_nacc_1843_update_completed__ps
      -- 
    ack_4473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1892_1843_buf_ack_1, ack => convolve_CP_4332_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_acc_var_1844_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_acc_var_1844_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_acc_var_1844_sample_start__ps
      -- CP-element group 54: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_acc_var_1844_sample_completed__ps
      -- 
    -- Element group convolve_CP_4332_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_acc_var_1844_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_acc_var_1844_update_start__ps
      -- 
    -- Element group convolve_CP_4332_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_acc_var_1844_update_completed__ps
      -- 
    convolve_CP_4332_elements(56) <= convolve_CP_4332_elements(57);
    -- CP-element group 57:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	56 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_acc_var_1844_update_completed_
      -- 
    -- Element group convolve_CP_4332_elements(57) is a control-delay.
    cp_element_57_delay: control_delay_element  generic map(name => " 57_delay", delay_value => 1)  port map(req => convolve_CP_4332_elements(55), ack => convolve_CP_4332_elements(57), clk => clk, reset =>reset);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	86 
    -- CP-element group 58: 	17 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	16 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_sample_start_
      -- 
    convolve_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(86) & convolve_CP_4332_elements(17);
      gj_convolve_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	14 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	88 
    -- CP-element group 59: 	91 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	18 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_update_start_
      -- 
    convolve_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(88) & convolve_CP_4332_elements(91);
      gj_convolve_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	17 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_sample_completed__ps
      -- 
    -- Element group convolve_CP_4332_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	87 
    -- CP-element group 61: 	90 
    -- CP-element group 61: 	19 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_update_completed__ps
      -- 
    -- Element group convolve_CP_4332_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	12 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_loopback_trigger
      -- 
    convolve_CP_4332_elements(62) <= convolve_CP_4332_elements(12);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_loopback_sample_req
      -- CP-element group 63: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_loopback_sample_req_ps
      -- 
    phi_stmt_1845_loopback_sample_req_4492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1845_loopback_sample_req_4492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(63), ack => phi_stmt_1845_req_1); -- 
    -- Element group convolve_CP_4332_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	13 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_entry_trigger
      -- 
    convolve_CP_4332_elements(64) <= convolve_CP_4332_elements(13);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_entry_sample_req
      -- CP-element group 65: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_entry_sample_req_ps
      -- 
    phi_stmt_1845_entry_sample_req_4495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1845_entry_sample_req_4495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(65), ack => phi_stmt_1845_req_0); -- 
    -- Element group convolve_CP_4332_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_phi_mux_ack
      -- CP-element group 66: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/phi_stmt_1845_phi_mux_ack_ps
      -- 
    phi_stmt_1845_phi_mux_ack_4498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1845_ack_0, ack => convolve_CP_4332_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1848_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1848_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1848_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1848_sample_completed_
      -- 
    -- Element group convolve_CP_4332_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1848_update_start__ps
      -- CP-element group 68: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1848_update_start_
      -- 
    -- Element group convolve_CP_4332_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1848_update_completed__ps
      -- 
    convolve_CP_4332_elements(69) <= convolve_CP_4332_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1848_update_completed_
      -- 
    -- Element group convolve_CP_4332_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convolve_CP_4332_elements(68), ack => convolve_CP_4332_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_sample_start__ps
      -- CP-element group 71: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_Sample/req
      -- 
    req_4519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(71), ack => n_out_count_1921_1849_buf_req_0); -- 
    -- Element group convolve_CP_4332_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_Update/req
      -- CP-element group 72: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_update_start__ps
      -- CP-element group 72: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_update_start_
      -- 
    req_4524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(72), ack => n_out_count_1921_1849_buf_req_1); -- 
    -- Element group convolve_CP_4332_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_sample_completed__ps
      -- CP-element group 73: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_sample_completed_
      -- 
    ack_4520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1921_1849_buf_ack_0, ack => convolve_CP_4332_elements(73)); -- 
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_update_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/R_n_out_count_1849_update_completed_
      -- 
    ack_4525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1921_1849_buf_ack_1, ack => convolve_CP_4332_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	78 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_Sample/rr
      -- 
    rr_4534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(75), ack => RPIPE_input_pipe1_1852_inst_req_0); -- 
    convolve_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(78);
      gj_convolve_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	17 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	95 
    -- CP-element group 76: 	99 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_update_start_
      -- CP-element group 76: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_Update/cr
      -- 
    cr_4539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(76), ack => RPIPE_input_pipe1_1852_inst_req_1); -- 
    convolve_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(77) & convolve_CP_4332_elements(17) & convolve_CP_4332_elements(95) & convolve_CP_4332_elements(99);
      gj_convolve_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	76 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_Sample/$exit
      -- 
    ra_4535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1852_inst_ack_0, ack => convolve_CP_4332_elements(77)); -- 
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	93 
    -- CP-element group 78: 	97 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: 	39 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_input_pipe1_1852_Update/ca
      -- 
    ca_4540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1852_inst_ack_1, ack => convolve_CP_4332_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	14 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_Sample/$entry
      -- 
    rr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(79), ack => RPIPE_kernel_pipe1_1859_inst_req_0); -- 
    convolve_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(82);
      gj_convolve_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	17 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	88 
    -- CP-element group 80: 	95 
    -- CP-element group 80: 	99 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_update_start_
      -- 
    cr_4553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(80), ack => RPIPE_kernel_pipe1_1859_inst_req_1); -- 
    convolve_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 15,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(81) & convolve_CP_4332_elements(17) & convolve_CP_4332_elements(88) & convolve_CP_4332_elements(95) & convolve_CP_4332_elements(99);
      gj_convolve_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	80 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_sample_completed_
      -- 
    ra_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1859_inst_ack_0, ack => convolve_CP_4332_elements(81)); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	87 
    -- CP-element group 82: 	93 
    -- CP-element group 82: 	97 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: 	39 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/RPIPE_kernel_pipe1_1859_Update/ca
      -- 
    ca_4554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1859_inst_ack_1, ack => convolve_CP_4332_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	14 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_Sample/rr
      -- 
    rr_4562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(83), ack => SUB_u32_u32_1873_inst_req_0); -- 
    convolve_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(14) & convolve_CP_4332_elements(85);
      gj_convolve_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	17 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	91 
    -- CP-element group 84: 	114 
    -- CP-element group 84: 	103 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_update_start_
      -- CP-element group 84: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_Update/cr
      -- 
    cr_4567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(84), ack => SUB_u32_u32_1873_inst_req_1); -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(17) & convolve_CP_4332_elements(91) & convolve_CP_4332_elements(114) & convolve_CP_4332_elements(103);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_Sample/ra
      -- 
    ra_4563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1873_inst_ack_0, ack => convolve_CP_4332_elements(85)); -- 
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	90 
    -- CP-element group 86: 	112 
    -- CP-element group 86: 	101 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	58 
    -- CP-element group 86: 	20 
    -- CP-element group 86: 	39 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/SUB_u32_u32_1873_Update/ca
      -- 
    ca_4568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1873_inst_ack_1, ack => convolve_CP_4332_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	82 
    -- CP-element group 87: 	61 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_Sample/$entry
      -- 
    req_4576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(87), ack => WPIPE_kernel_pipe1_1907_inst_req_0); -- 
    convolve_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(82) & convolve_CP_4332_elements(61) & convolve_CP_4332_elements(89);
      gj_convolve_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	80 
    -- CP-element group 88: 	59 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_Sample/ack
      -- CP-element group 88: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_Sample/$exit
      -- 
    ack_4577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1907_inst_ack_0, ack => convolve_CP_4332_elements(88)); -- 
    req_4581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(88), ack => WPIPE_kernel_pipe1_1907_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	124 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_Update/ack
      -- CP-element group 89: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_kernel_pipe1_1907_update_completed_
      -- 
    ack_4582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1907_inst_ack_1, ack => convolve_CP_4332_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	86 
    -- CP-element group 90: 	61 
    -- CP-element group 90: 	25 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_Sample/req
      -- 
    req_4590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(90), ack => WPIPE_input_done_pipe_1928_inst_req_0); -- 
    convolve_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(86) & convolve_CP_4332_elements(61) & convolve_CP_4332_elements(25) & convolve_CP_4332_elements(92);
      gj_convolve_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	84 
    -- CP-element group 91: 	59 
    -- CP-element group 91: 	21 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_Update/req
      -- 
    ack_4591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1928_inst_ack_0, ack => convolve_CP_4332_elements(91)); -- 
    req_4595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(91), ack => WPIPE_input_done_pipe_1928_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	124 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_Update/ack
      -- CP-element group 92: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_input_done_pipe_1928_update_completed_
      -- 
    ack_4596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1928_inst_ack_1, ack => convolve_CP_4332_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	78 
    -- CP-element group 93: 	82 
    -- CP-element group 93: 	44 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_Sample/rr
      -- 
    rr_4604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(93), ack => slice_1933_inst_req_0); -- 
    convolve_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(78) & convolve_CP_4332_elements(82) & convolve_CP_4332_elements(44) & convolve_CP_4332_elements(95);
      gj_convolve_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	107 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_Update/cr
      -- 
    cr_4609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(94), ack => slice_1933_inst_req_1); -- 
    convolve_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4332_elements(107);
      gj_convolve_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	76 
    -- CP-element group 95: 	80 
    -- CP-element group 95: 	40 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_Sample/ra
      -- 
    ra_4605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1933_inst_ack_0, ack => convolve_CP_4332_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	105 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1933_Update/ca
      -- 
    ca_4610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1933_inst_ack_1, ack => convolve_CP_4332_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	78 
    -- CP-element group 97: 	82 
    -- CP-element group 97: 	44 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_Sample/rr
      -- 
    rr_4618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(97), ack => slice_1937_inst_req_0); -- 
    convolve_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(78) & convolve_CP_4332_elements(82) & convolve_CP_4332_elements(44) & convolve_CP_4332_elements(99);
      gj_convolve_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	118 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_Update/$entry
      -- 
    cr_4623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(98), ack => slice_1937_inst_req_1); -- 
    convolve_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4332_elements(118);
      gj_convolve_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	76 
    -- CP-element group 99: 	80 
    -- CP-element group 99: 	40 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_Sample/$exit
      -- 
    ra_4619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1937_inst_ack_0, ack => convolve_CP_4332_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	116 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/slice_1937_Update/$exit
      -- 
    ca_4624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1937_inst_ack_1, ack => convolve_CP_4332_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	86 
    -- CP-element group 101: 	25 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_Sample/req
      -- CP-element group 101: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_sample_start_
      -- 
    req_4632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(101), ack => W_next_sum_1915_delayed_1_0_1939_inst_req_0); -- 
    convolve_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(86) & convolve_CP_4332_elements(25) & convolve_CP_4332_elements(103);
      gj_convolve_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	107 
    -- CP-element group 102: 	110 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_Update/req
      -- 
    req_4637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(102), ack => W_next_sum_1915_delayed_1_0_1939_inst_req_1); -- 
    convolve_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(107) & convolve_CP_4332_elements(110);
      gj_convolve_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	84 
    -- CP-element group 103: 	21 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_Sample/ack
      -- 
    ack_4633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1915_delayed_1_0_1939_inst_ack_0, ack => convolve_CP_4332_elements(103)); -- 
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	109 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1941_Update/ack
      -- 
    ack_4638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1915_delayed_1_0_1939_inst_ack_1, ack => convolve_CP_4332_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	96 
    -- CP-element group 105: 	104 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_sample_start_
      -- 
    rr_4646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(105), ack => type_cast_1945_inst_req_0); -- 
    convolve_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(96) & convolve_CP_4332_elements(104) & convolve_CP_4332_elements(107);
      gj_convolve_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	110 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_update_start_
      -- CP-element group 106: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_Update/cr
      -- 
    cr_4651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(106), ack => type_cast_1945_inst_req_1); -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4332_elements(110);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	94 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_sample_completed_
      -- 
    ra_4647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_0, ack => convolve_CP_4332_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1945_update_completed_
      -- 
    ca_4652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_1, ack => convolve_CP_4332_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: 	104 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	122 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_Sample/req
      -- CP-element group 109: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_Sample/$entry
      -- 
    req_4660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(109), ack => WPIPE_maxpool_output_pipe_1943_inst_req_0); -- 
    convolve_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(108) & convolve_CP_4332_elements(104) & convolve_CP_4332_elements(122);
      gj_convolve_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	102 
    -- CP-element group 110: 	106 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_Sample/ack
      -- CP-element group 110: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_Update/req
      -- 
    ack_4661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1943_inst_ack_0, ack => convolve_CP_4332_elements(110)); -- 
    req_4665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(110), ack => WPIPE_maxpool_output_pipe_1943_inst_req_1); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	120 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1943_Update/ack
      -- 
    ack_4666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1943_inst_ack_1, ack => convolve_CP_4332_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	86 
    -- CP-element group 112: 	25 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_Sample/req
      -- 
    req_4674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(112), ack => W_next_sum_1920_delayed_1_0_1947_inst_req_0); -- 
    convolve_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(86) & convolve_CP_4332_elements(25) & convolve_CP_4332_elements(114);
      gj_convolve_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	118 
    -- CP-element group 113: 	121 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_Update/req
      -- 
    req_4679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(113), ack => W_next_sum_1920_delayed_1_0_1947_inst_req_1); -- 
    convolve_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(118) & convolve_CP_4332_elements(121);
      gj_convolve_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	84 
    -- CP-element group 114: 	21 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_Sample/ack
      -- 
    ack_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1920_delayed_1_0_1947_inst_ack_0, ack => convolve_CP_4332_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	120 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/assign_stmt_1949_Update/ack
      -- 
    ack_4680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1920_delayed_1_0_1947_inst_ack_1, ack => convolve_CP_4332_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: 	100 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_Sample/rr
      -- 
    rr_4688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(116), ack => type_cast_1953_inst_req_0); -- 
    convolve_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(115) & convolve_CP_4332_elements(100) & convolve_CP_4332_elements(118);
      gj_convolve_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_update_start_
      -- CP-element group 117: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_Update/cr
      -- 
    cr_4693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(117), ack => type_cast_1953_inst_req_1); -- 
    convolve_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4332_elements(121);
      gj_convolve_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	98 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_Sample/ra
      -- 
    ra_4689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_0, ack => convolve_CP_4332_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/type_cast_1953_Update/ca
      -- 
    ca_4694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_1, ack => convolve_CP_4332_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	111 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	119 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_Sample/req
      -- 
    req_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(120), ack => WPIPE_maxpool_output_pipe_1951_inst_req_0); -- 
    convolve_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(111) & convolve_CP_4332_elements(115) & convolve_CP_4332_elements(119) & convolve_CP_4332_elements(122);
      gj_convolve_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	113 
    -- CP-element group 121: 	117 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_update_start_
      -- CP-element group 121: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_Sample/ack
      -- CP-element group 121: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_Update/req
      -- 
    ack_4703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1951_inst_ack_0, ack => convolve_CP_4332_elements(121)); -- 
    req_4707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4332_elements(121), ack => WPIPE_maxpool_output_pipe_1951_inst_req_1); -- 
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	109 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/WPIPE_maxpool_output_pipe_1951_Update/ack
      -- 
    ack_4708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1951_inst_ack_1, ack => convolve_CP_4332_elements(122)); -- 
    -- CP-element group 123:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	14 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	15 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_4332_elements(123) is a control-delay.
    cp_element_123_delay: control_delay_element  generic map(name => " 123_delay", delay_value => 1)  port map(req => convolve_CP_4332_elements(14), ack => convolve_CP_4332_elements(123), clk => clk, reset =>reset);
    -- CP-element group 124:  join  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	89 
    -- CP-element group 124: 	92 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	11 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1819/do_while_stmt_1835/do_while_stmt_1835_loop_body/$exit
      -- 
    convolve_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4332_elements(89) & convolve_CP_4332_elements(92) & convolve_CP_4332_elements(122);
      gj_convolve_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4332_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	10 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1819/do_while_stmt_1835/loop_exit/$exit
      -- CP-element group 125: 	 branch_block_stmt_1819/do_while_stmt_1835/loop_exit/ack
      -- 
    ack_4713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1835_branch_ack_0, ack => convolve_CP_4332_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	10 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1819/do_while_stmt_1835/loop_taken/$exit
      -- CP-element group 126: 	 branch_block_stmt_1819/do_while_stmt_1835/loop_taken/ack
      -- 
    ack_4717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1835_branch_ack_1, ack => convolve_CP_4332_elements(126)); -- 
    -- CP-element group 127:  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	8 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1819/do_while_stmt_1835/$exit
      -- 
    convolve_CP_4332_elements(127) <= convolve_CP_4332_elements(8);
    convolve_do_while_stmt_1835_terminator_4718: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1835_terminator_4718", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_4332_elements(11),loop_continue => convolve_CP_4332_elements(126),loop_terminate => convolve_CP_4332_elements(125),loop_back => convolve_CP_4332_elements(9),loop_exit => convolve_CP_4332_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1837_phi_seq_4438_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4332_elements(26);
      convolve_CP_4332_elements(31)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4332_elements(33);
      convolve_CP_4332_elements(32)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4332_elements(34);
      convolve_CP_4332_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4332_elements(28);
      convolve_CP_4332_elements(35)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4332_elements(35);
      convolve_CP_4332_elements(36)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4332_elements(37);
      convolve_CP_4332_elements(29) <= phi_mux_reqs(1);
      phi_stmt_1837_phi_seq_4438 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1837_phi_seq_4438") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4332_elements(22), 
          phi_sample_ack => convolve_CP_4332_elements(23), 
          phi_update_req => convolve_CP_4332_elements(24), 
          phi_update_ack => convolve_CP_4332_elements(25), 
          phi_mux_ack => convolve_CP_4332_elements(30), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1841_phi_seq_4482_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4332_elements(45);
      convolve_CP_4332_elements(50)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4332_elements(52);
      convolve_CP_4332_elements(51)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4332_elements(53);
      convolve_CP_4332_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4332_elements(47);
      convolve_CP_4332_elements(54)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4332_elements(54);
      convolve_CP_4332_elements(55)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4332_elements(56);
      convolve_CP_4332_elements(48) <= phi_mux_reqs(1);
      phi_stmt_1841_phi_seq_4482 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1841_phi_seq_4482") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4332_elements(41), 
          phi_sample_ack => convolve_CP_4332_elements(42), 
          phi_update_req => convolve_CP_4332_elements(43), 
          phi_update_ack => convolve_CP_4332_elements(44), 
          phi_mux_ack => convolve_CP_4332_elements(49), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1845_phi_seq_4526_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4332_elements(64);
      convolve_CP_4332_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4332_elements(67);
      convolve_CP_4332_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4332_elements(69);
      convolve_CP_4332_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4332_elements(62);
      convolve_CP_4332_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4332_elements(73);
      convolve_CP_4332_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4332_elements(74);
      convolve_CP_4332_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1845_phi_seq_4526 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1845_phi_seq_4526") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4332_elements(16), 
          phi_sample_ack => convolve_CP_4332_elements(60), 
          phi_update_req => convolve_CP_4332_elements(18), 
          phi_update_ack => convolve_CP_4332_elements(61), 
          phi_mux_ack => convolve_CP_4332_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4390_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_4332_elements(12);
        preds(1)  <= convolve_CP_4332_elements(13);
        entry_tmerge_4390 : transition_merge -- 
          generic map(name => " entry_tmerge_4390")
          port map (preds => preds, symbol_out => convolve_CP_4332_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1917_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_1898_wire : std_logic_vector(31 downto 0);
    signal MUX_1918_wire : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_1853_1853_delayed_1_0_1874 : std_logic_vector(31 downto 0);
    signal acc_1841 : std_logic_vector(15 downto 0);
    signal acc_val_1886 : std_logic_vector(15 downto 0);
    signal acc_val_dn_1938 : std_logic_vector(7 downto 0);
    signal acc_val_up_1934 : std_logic_vector(7 downto 0);
    signal acc_var_1834 : std_logic_vector(15 downto 0);
    signal all_done_flag_1926 : std_logic_vector(0 downto 0);
    signal iread_1853 : std_logic_vector(15 downto 0);
    signal ival_1857 : std_logic_vector(15 downto 0);
    signal konst_1872_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1889_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1895_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1897_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1916_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1929_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1956_wire_constant : std_logic_vector(0 downto 0);
    signal kread_1860 : std_logic_vector(15 downto 0);
    signal kval_1864 : std_logic_vector(15 downto 0);
    signal mcount_var_1829 : std_logic_vector(31 downto 0);
    signal mul_val_1869 : std_logic_vector(15 downto 0);
    signal mycount_1837 : std_logic_vector(31 downto 0);
    signal n_out_count_1921 : std_logic_vector(15 downto 0);
    signal n_out_count_1921_1849_buffered : std_logic_vector(15 downto 0);
    signal nacc_1892 : std_logic_vector(15 downto 0);
    signal nacc_1892_1843_buffered : std_logic_vector(15 downto 0);
    signal next_sum_1879 : std_logic_vector(0 downto 0);
    signal next_sum_1915_delayed_1_0_1941 : std_logic_vector(0 downto 0);
    signal next_sum_1920_delayed_1_0_1949 : std_logic_vector(0 downto 0);
    signal nmycount_1900 : std_logic_vector(31 downto 0);
    signal nmycount_1900_1839_buffered : std_logic_vector(31 downto 0);
    signal num_out_1822 : std_logic_vector(15 downto 0);
    signal out_count_1845 : std_logic_vector(15 downto 0);
    signal out_done_flag_1905 : std_logic_vector(0 downto 0);
    signal size_1825 : std_logic_vector(31 downto 0);
    signal type_cast_1848_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1882_wire : std_logic_vector(15 downto 0);
    signal type_cast_1884_wire : std_logic_vector(15 downto 0);
    signal type_cast_1914_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1945_wire : std_logic_vector(7 downto 0);
    signal type_cast_1953_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    acc_var_1834 <= "0000000000000000";
    konst_1872_wire_constant <= "00000000000000000000000000000001";
    konst_1889_wire_constant <= "0000000000000000";
    konst_1895_wire_constant <= "00000000000000000000000000000000";
    konst_1897_wire_constant <= "00000000000000000000000000000001";
    konst_1916_wire_constant <= "0000000000000001";
    konst_1929_wire_constant <= "1";
    konst_1956_wire_constant <= "1";
    mcount_var_1829 <= "00000000000000000000000000000000";
    type_cast_1848_wire_constant <= "0000000000000001";
    type_cast_1914_wire_constant <= "0000000000000001";
    phi_stmt_1837: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_1900_1839_buffered & mcount_var_1829;
      req <= phi_stmt_1837_req_0 & phi_stmt_1837_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1837",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1837_ack_0,
          idata => idata,
          odata => mycount_1837,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1837
    phi_stmt_1841: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nacc_1892_1843_buffered & acc_var_1834;
      req <= phi_stmt_1841_req_0 & phi_stmt_1841_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1841",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1841_ack_0,
          idata => idata,
          odata => acc_1841,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1841
    phi_stmt_1845: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1848_wire_constant & n_out_count_1921_1849_buffered;
      req <= phi_stmt_1845_req_0 & phi_stmt_1845_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1845",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1845_ack_0,
          idata => idata,
          odata => out_count_1845,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1845
    -- flow-through select operator MUX_1891_inst
    nacc_1892 <= konst_1889_wire_constant when (next_sum_1879(0) /=  '0') else acc_val_1886;
    -- flow-through select operator MUX_1899_inst
    nmycount_1900 <= konst_1895_wire_constant when (next_sum_1879(0) /=  '0') else ADD_u32_u32_1898_wire;
    -- flow-through select operator MUX_1918_inst
    MUX_1918_wire <= type_cast_1914_wire_constant when (out_done_flag_1905(0) /=  '0') else ADD_u16_u16_1917_wire;
    -- flow-through select operator MUX_1920_inst
    n_out_count_1921 <= MUX_1918_wire when (next_sum_1879(0) /=  '0') else out_count_1845;
    slice_1933_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1933_inst_req_0;
      slice_1933_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1933_inst_req_1;
      slice_1933_inst_ack_1<= update_ack(0);
      slice_1933_inst: SliceSplitProtocol generic map(name => "slice_1933_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1886, dout => acc_val_up_1934, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1937_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1937_inst_req_0;
      slice_1937_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1937_inst_req_1;
      slice_1937_inst_ack_1<= update_ack(0);
      slice_1937_inst: SliceSplitProtocol generic map(name => "slice_1937_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1886, dout => acc_val_dn_1938, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_next_sum_1915_delayed_1_0_1939_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1915_delayed_1_0_1939_inst_req_0;
      W_next_sum_1915_delayed_1_0_1939_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1915_delayed_1_0_1939_inst_req_1;
      W_next_sum_1915_delayed_1_0_1939_inst_ack_1<= rack(0);
      W_next_sum_1915_delayed_1_0_1939_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1915_delayed_1_0_1939_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1879,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1915_delayed_1_0_1941,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_next_sum_1920_delayed_1_0_1947_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1920_delayed_1_0_1947_inst_req_0;
      W_next_sum_1920_delayed_1_0_1947_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1920_delayed_1_0_1947_inst_req_1;
      W_next_sum_1920_delayed_1_0_1947_inst_ack_1<= rack(0);
      W_next_sum_1920_delayed_1_0_1947_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1920_delayed_1_0_1947_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1879,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1920_delayed_1_0_1949,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_out_count_1921_1849_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_out_count_1921_1849_buf_req_0;
      n_out_count_1921_1849_buf_ack_0<= wack(0);
      rreq(0) <= n_out_count_1921_1849_buf_req_1;
      n_out_count_1921_1849_buf_ack_1<= rack(0);
      n_out_count_1921_1849_buf : InterlockBuffer generic map ( -- 
        name => "n_out_count_1921_1849_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_out_count_1921,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_out_count_1921_1849_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_1892_1843_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_1892_1843_buf_req_0;
      nacc_1892_1843_buf_ack_0<= wack(0);
      rreq(0) <= nacc_1892_1843_buf_req_1;
      nacc_1892_1843_buf_ack_1<= rack(0);
      nacc_1892_1843_buf : InterlockBuffer generic map ( -- 
        name => "nacc_1892_1843_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_1892,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_1892_1843_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_1900_1839_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_1900_1839_buf_req_0;
      nmycount_1900_1839_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_1900_1839_buf_req_1;
      nmycount_1900_1839_buf_ack_1<= rack(0);
      nmycount_1900_1839_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_1900_1839_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_1900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_1900_1839_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1856_inst
    process(iread_1853) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread_1853(15 downto 0);
      ival_1857 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1863_inst
    process(kread_1860) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread_1860(15 downto 0);
      kval_1864 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1882_inst
    process(acc_1841) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := acc_1841(15 downto 0);
      type_cast_1882_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1884_inst
    process(mul_val_1869) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mul_val_1869(15 downto 0);
      type_cast_1884_wire <= tmp_var; -- 
    end process;
    type_cast_1945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1945_inst_req_0;
      type_cast_1945_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1945_inst_req_1;
      type_cast_1945_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1915_delayed_1_0_1941(0);
      type_cast_1945_inst_gI: SplitGuardInterface generic map(name => "type_cast_1945_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_up_1934,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1945_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1953_inst_req_0;
      type_cast_1953_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1953_inst_req_1;
      type_cast_1953_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1920_delayed_1_0_1949(0);
      type_cast_1953_inst_gI: SplitGuardInterface generic map(name => "type_cast_1953_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1953_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1953_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_dn_1938,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1953_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1835_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1956_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1835_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1835_branch_req_0,
          ack0 => do_while_stmt_1835_branch_ack_0,
          ack1 => do_while_stmt_1835_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_1885_inst
    process(type_cast_1882_wire, type_cast_1884_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_1882_wire, type_cast_1884_wire, tmp_var);
      acc_val_1886 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1917_inst
    process(out_count_1845) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_count_1845, konst_1916_wire_constant, tmp_var);
      ADD_u16_u16_1917_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1898_inst
    process(mycount_1837) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_1837, konst_1897_wire_constant, tmp_var);
      ADD_u32_u32_1898_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1925_inst
    process(out_done_flag_1905, next_sum_1879) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_1905, next_sum_1879, tmp_var);
      all_done_flag_1926 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1904_inst
    process(out_count_1845, num_out_1822) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(out_count_1845, num_out_1822, tmp_var);
      out_done_flag_1905 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1878_inst
    process(mycount_1837, SUB_u32_u32_1853_1853_delayed_1_0_1874) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycount_1837, SUB_u32_u32_1853_1853_delayed_1_0_1874, tmp_var);
      next_sum_1879 <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_1868_inst
    process(kval_1864, ival_1857) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval_1864, ival_1857, tmp_var);
      mul_val_1869 <= tmp_var; --
    end process;
    -- shared split operator group (7) : SUB_u32_u32_1873_inst 
    ApIntSub_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= size_1825;
      SUB_u32_u32_1853_1853_delayed_1_0_1874 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_1873_inst_req_0;
      SUB_u32_u32_1873_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_1873_inst_req_1;
      SUB_u32_u32_1873_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_7_gI: SplitGuardInterface generic map(name => "ApIntSub_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared inport operator group (0) : RPIPE_input_pipe1_1852_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1852_inst_req_0;
      RPIPE_input_pipe1_1852_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1852_inst_req_1;
      RPIPE_input_pipe1_1852_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iread_1853 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_kernel_pipe1_1859_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_1859_inst_req_0;
      RPIPE_kernel_pipe1_1859_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_1859_inst_req_1;
      RPIPE_kernel_pipe1_1859_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      kread_1860 <= data_out(15 downto 0);
      kernel_pipe1_read_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_num_out_pipe_1821_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1821_inst_req_0;
      RPIPE_num_out_pipe_1821_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1821_inst_req_1;
      RPIPE_num_out_pipe_1821_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      num_out_1822 <= data_out(15 downto 0);
      num_out_pipe_read_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_2: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_size_pipe_1824_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1824_inst_req_0;
      RPIPE_size_pipe_1824_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1824_inst_req_1;
      RPIPE_size_pipe_1824_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      size_1825 <= data_out(31 downto 0);
      size_pipe_read_3_gI: SplitGuardInterface generic map(name => "size_pipe_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_3: InputPortRevised -- 
        generic map ( name => "size_pipe_read_3", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_input_done_pipe_1928_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_1928_inst_req_0;
      WPIPE_input_done_pipe_1928_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_1928_inst_req_1;
      WPIPE_input_done_pipe_1928_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= all_done_flag_1926(0);
      data_in <= konst_1929_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe1_1907_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_1907_inst_req_0;
      WPIPE_kernel_pipe1_1907_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_1907_inst_req_1;
      WPIPE_kernel_pipe1_1907_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not out_done_flag_1905(0);
      data_in <= kread_1860;
      kernel_pipe1_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_maxpool_output_pipe_1943_inst WPIPE_maxpool_output_pipe_1951_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1943_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1951_inst_req_0;
      WPIPE_maxpool_output_pipe_1943_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1951_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1943_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1951_inst_req_1;
      WPIPE_maxpool_output_pipe_1943_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1951_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= next_sum_1920_delayed_1_0_1949(0);
      guard_vector(1)  <= next_sum_1915_delayed_1_0_1941(0);
      data_in <= type_cast_1945_wire & type_cast_1953_wire;
      maxpool_output_pipe_write_2_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    end_add : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 128)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal end_add_buffer :  std_logic_vector(63 downto 0);
  signal end_add_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_676_start: Boolean;
  signal loadKernelChannel_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal addr_of_398_final_reg_req_0 : boolean;
  signal phi_stmt_356_req_1 : boolean;
  signal type_cast_432_inst_ack_0 : boolean;
  signal do_while_stmt_350_branch_ack_0 : boolean;
  signal my_fetch_339_359_buf_req_1 : boolean;
  signal nfetch_val_419_358_buf_req_0 : boolean;
  signal addr_of_398_final_reg_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_req_0 : boolean;
  signal array_obj_ref_397_index_offset_req_0 : boolean;
  signal WPIPE_size_pipe_428_inst_ack_0 : boolean;
  signal do_while_stmt_350_branch_ack_1 : boolean;
  signal addr_of_398_final_reg_req_1 : boolean;
  signal type_cast_432_inst_req_0 : boolean;
  signal WPIPE_size_pipe_428_inst_req_1 : boolean;
  signal addr_of_398_final_reg_ack_1 : boolean;
  signal WPIPE_size_pipe_428_inst_ack_1 : boolean;
  signal my_fetch_339_359_buf_ack_0 : boolean;
  signal phi_stmt_356_ack_0 : boolean;
  signal array_obj_ref_397_index_offset_ack_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_req_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_ack_0 : boolean;
  signal nfetch_val_419_358_buf_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_ack_1 : boolean;
  signal phi_stmt_356_req_0 : boolean;
  signal ptr_deref_406_load_0_req_0 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_req_0 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_ack_0 : boolean;
  signal nfetch_val_419_358_buf_req_1 : boolean;
  signal my_fetch_339_359_buf_ack_1 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_req_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_req_1 : boolean;
  signal array_obj_ref_397_index_offset_req_1 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_req_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_ack_1 : boolean;
  signal array_obj_ref_397_index_offset_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_ack_0 : boolean;
  signal my_fetch_339_359_buf_req_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_ack_1 : boolean;
  signal ptr_deref_406_load_0_ack_0 : boolean;
  signal nfetch_val_419_358_buf_ack_1 : boolean;
  signal type_cast_432_inst_req_1 : boolean;
  signal WPIPE_size_pipe_428_inst_req_0 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_ack_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_req_1 : boolean;
  signal array_obj_ref_333_index_offset_req_0 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_ack_0 : boolean;
  signal array_obj_ref_333_index_offset_ack_0 : boolean;
  signal array_obj_ref_333_index_offset_req_1 : boolean;
  signal array_obj_ref_333_index_offset_ack_1 : boolean;
  signal type_cast_432_inst_ack_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_req_0 : boolean;
  signal addr_of_334_final_reg_req_0 : boolean;
  signal addr_of_334_final_reg_ack_0 : boolean;
  signal addr_of_334_final_reg_req_1 : boolean;
  signal addr_of_334_final_reg_ack_1 : boolean;
  signal ptr_deref_406_load_0_ack_1 : boolean;
  signal ptr_deref_406_load_0_req_1 : boolean;
  signal ptr_deref_338_load_0_req_0 : boolean;
  signal ptr_deref_338_load_0_ack_0 : boolean;
  signal start_add_355_buf_ack_1 : boolean;
  signal ptr_deref_338_load_0_req_1 : boolean;
  signal ptr_deref_338_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_347_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_347_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_347_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_347_inst_ack_1 : boolean;
  signal do_while_stmt_350_branch_req_0 : boolean;
  signal phi_stmt_352_req_0 : boolean;
  signal phi_stmt_352_req_1 : boolean;
  signal phi_stmt_352_ack_0 : boolean;
  signal nmycount_374_354_buf_req_0 : boolean;
  signal nmycount_374_354_buf_ack_0 : boolean;
  signal nmycount_374_354_buf_req_1 : boolean;
  signal nmycount_374_354_buf_ack_1 : boolean;
  signal start_add_355_buf_req_0 : boolean;
  signal start_add_355_buf_ack_0 : boolean;
  signal start_add_355_buf_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 128) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= end_add;
  end_add_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(tag_length + 127 downto 128) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 127 downto 128);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_676: Block -- control-path 
    signal loadKernelChannel_CP_676_elements: BooleanArray(94 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_676_elements(0) <= loadKernelChannel_CP_676_start;
    loadKernelChannel_CP_676_symbol <= loadKernelChannel_CP_676_elements(94);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_update_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resized_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_computed_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_update_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_sample_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/rr
      -- 
    rr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => RPIPE_input_done_pipe_347_inst_req_0); -- 
    req_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_333_index_offset_req_1); -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_333_index_offset_req_0); -- 
    req_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => addr_of_334_final_reg_req_1); -- 
    cr_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => ptr_deref_338_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/ack
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_333_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_sample_start_
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_offset_calculated
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/$entry
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/req
      -- 
    ack_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_333_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(2)); -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(2), ack => addr_of_334_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_sample_completed_
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/$exit
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/ack
      -- 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_334_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_update_completed_
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_sample_start_
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_address_resized
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/rr
      -- 
    ack_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_334_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(4)); -- 
    rr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(4), ack => ptr_deref_338_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_sample_completed_
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/ra
      -- 
    ra_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_338_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_update_completed_
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/merge_ack
      -- 
    ca_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_338_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_sample_completed_
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_update_start_
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/ra
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/$entry
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/cr
      -- 
    ra_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_347_inst_ack_0, ack => loadKernelChannel_CP_676_elements(7)); -- 
    cr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(7), ack => RPIPE_input_done_pipe_347_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_update_completed_
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/$exit
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/ca
      -- 
    ca_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_347_inst_ack_1, ack => loadKernelChannel_CP_676_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_328_to_assign_stmt_348/$exit
      -- CP-element group 9: 	 branch_block_stmt_349/$entry
      -- CP-element group 9: 	 branch_block_stmt_349/branch_block_stmt_349__entry__
      -- CP-element group 9: 	 branch_block_stmt_349/do_while_stmt_350__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(6) & loadKernelChannel_CP_676_elements(1) & loadKernelChannel_CP_676_elements(8);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	90 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	91 
    -- CP-element group 10: 	92 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Sample/rr
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Update/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_update_start_
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_sample_start_
      -- CP-element group 10: 	 assign_stmt_433/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_349/$exit
      -- CP-element group 10: 	 branch_block_stmt_349/branch_block_stmt_349__exit__
      -- CP-element group 10: 	 branch_block_stmt_349/do_while_stmt_350__exit__
      -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_432_inst_req_0); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_432_inst_req_1); -- 
    loadKernelChannel_CP_676_elements(10) <= loadKernelChannel_CP_676_elements(90);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_349/do_while_stmt_350/$entry
      -- CP-element group 11: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350__entry__
      -- 
    loadKernelChannel_CP_676_elements(11) <= loadKernelChannel_CP_676_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	90 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350__exit__
      -- 
    -- Element group loadKernelChannel_CP_676_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_349/do_while_stmt_350/loop_back
      -- 
    -- Element group loadKernelChannel_CP_676_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	88 
    -- CP-element group 14: 	89 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/$entry
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/condition_done
      -- 
    loadKernelChannel_CP_676_elements(14) <= loadKernelChannel_CP_676_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	87 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_349/do_while_stmt_350/loop_body_done
      -- 
    loadKernelChannel_CP_676_elements(15) <= loadKernelChannel_CP_676_elements(87);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_676_elements(16) <= loadKernelChannel_CP_676_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	31 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_676_elements(17) <= loadKernelChannel_CP_676_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	43 
    -- CP-element group 18: 	86 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	64 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_676_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	86 
    -- CP-element group 19: 	28 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/condition_evaluated
      -- 
    condition_evaluated_813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(19), ack => do_while_stmt_350_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(23) & loadKernelChannel_CP_676_elements(86) & loadKernelChannel_CP_676_elements(28);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	42 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	26 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_start__ps
      -- CP-element group 20: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_sample_req
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(24) & loadKernelChannel_CP_676_elements(42) & loadKernelChannel_CP_676_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	27 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	75 
    -- CP-element group 21: 	79 
    -- CP-element group 21: 	87 
    -- CP-element group 21: 	83 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	42 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(27) & loadKernelChannel_CP_676_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	43 
    -- CP-element group 22: 	25 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_update_req
      -- CP-element group 22: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_start__ps
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(43) & loadKernelChannel_CP_676_elements(25);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(28) & loadKernelChannel_CP_676_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	66 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	80 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(28) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(72) & loadKernelChannel_CP_676_elements(80);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	20 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_start__ps
      -- 
    loadKernelChannel_CP_676_elements(26) <= loadKernelChannel_CP_676_elements(20);
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	21 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	19 
    -- CP-element group 28: 	23 
    -- CP-element group 28: 	78 
    -- CP-element group 28: 	60 
    -- CP-element group 28: 	66 
    -- CP-element group 28: 	70 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (15) 
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/scale_rename_req
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/$entry
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/index_resize_ack
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/scale_rename_ack
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/index_resize_req
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/$exit
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/$exit
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/$entry
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_computed_1
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scaled_1
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resized_1
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_completed__ps
      -- 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(28), ack => array_obj_ref_397_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	16 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_trigger
      -- 
    loadKernelChannel_CP_676_elements(29) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 30:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_sample_req
      -- CP-element group 30: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_sample_req_ps
      -- 
    phi_stmt_352_loopback_sample_req_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_352_loopback_sample_req_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(30), ack => phi_stmt_352_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(30) is bound as output of CP function.
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	17 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_trigger
      -- 
    loadKernelChannel_CP_676_elements(31) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 32:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_sample_req
      -- CP-element group 32: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_sample_req_ps
      -- 
    phi_stmt_352_entry_sample_req_831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_352_entry_sample_req_831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(32), ack => phi_stmt_352_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_phi_mux_ack
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_phi_mux_ack_ps
      -- 
    phi_stmt_352_phi_mux_ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_352_ack_0, ack => loadKernelChannel_CP_676_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/req
      -- 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(34), ack => nmycount_374_354_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_start_
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/req
      -- 
    req_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(35), ack => nmycount_374_354_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/ack
      -- 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_374_354_buf_ack_0, ack => loadKernelChannel_CP_676_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/ack
      -- 
    ack_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_374_354_buf_ack_1, ack => loadKernelChannel_CP_676_elements(37)); -- 
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_start__ps
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/req
      -- 
    req_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(38), ack => start_add_355_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_start__ps
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_start_
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/req
      -- 
    req_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(39), ack => start_add_355_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/ack
      -- 
    ack_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_355_buf_ack_0, ack => loadKernelChannel_CP_676_elements(40)); -- 
    -- CP-element group 41:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/$exit
      -- 
    ack_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_355_buf_ack_1, ack => loadKernelChannel_CP_676_elements(41)); -- 
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	21 
    -- CP-element group 42: 	77 
    -- CP-element group 42: 	81 
    -- CP-element group 42: 	85 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	20 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	18 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	61 
    -- CP-element group 43: 	84 
    -- CP-element group 43: 	46 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	22 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_start_
      -- 
    loadKernelChannel_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(84) & loadKernelChannel_CP_676_elements(46);
      gj_loadKernelChannel_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_start__ps
      -- 
    loadKernelChannel_CP_676_elements(45) <= loadKernelChannel_CP_676_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	82 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	43 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_completed_
      -- 
    -- Element group loadKernelChannel_CP_676_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_trigger
      -- 
    loadKernelChannel_CP_676_elements(47) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_sample_req_ps
      -- CP-element group 48: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_sample_req
      -- 
    phi_stmt_356_loopback_sample_req_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_356_loopback_sample_req_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(48), ack => phi_stmt_356_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_trigger
      -- 
    loadKernelChannel_CP_676_elements(49) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_sample_req_ps
      -- 
    phi_stmt_356_entry_sample_req_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_356_entry_sample_req_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(50), ack => phi_stmt_356_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_phi_mux_ack_ps
      -- 
    phi_stmt_356_phi_mux_ack_888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_356_ack_0, ack => loadKernelChannel_CP_676_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/$entry
      -- 
    req_901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(52), ack => nfetch_val_419_358_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_start_
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/req
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/$entry
      -- 
    req_906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(53), ack => nfetch_val_419_358_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_completed_
      -- 
    ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_419_358_buf_ack_0, ack => loadKernelChannel_CP_676_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/ack
      -- 
    ack_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_419_358_buf_ack_1, ack => loadKernelChannel_CP_676_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_start_
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(56), ack => my_fetch_339_359_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/req
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_start_
      -- 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(57), ack => my_fetch_339_359_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_completed_
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_339_359_buf_ack_0, ack => loadKernelChannel_CP_676_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_completed__ps
      -- 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_339_359_buf_ack_1, ack => loadKernelChannel_CP_676_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	28 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_sample_start_
      -- 
    req_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(60), ack => WPIPE_kernel_pipe1_381_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(28) & loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	43 
    -- CP-element group 61: 	25 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/req
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_update_start_
      -- 
    ack_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_381_inst_ack_0, ack => loadKernelChannel_CP_676_elements(61)); -- 
    req_939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(61), ack => WPIPE_kernel_pipe1_381_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	87 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/ack
      -- 
    ack_940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_381_inst_ack_1, ack => loadKernelChannel_CP_676_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	67 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	68 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/req
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/$entry
      -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(63), ack => addr_of_398_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	18 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	76 
    -- CP-element group 64: 	69 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/req
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_update_start_
      -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(64), ack => addr_of_398_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(76) & loadKernelChannel_CP_676_elements(69);
      gj_loadKernelChannel_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_update_start
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/req
      -- 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(65), ack => array_obj_ref_397_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	25 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_sample_complete
      -- 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_397_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	63 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (8) 
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/sum_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/$entry
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/$exit
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/sum_rename_req
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_offset_calculated
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_root_address_calculated
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_397_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	63 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/$exit
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/ack
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_sample_completed_
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_398_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	64 
    -- CP-element group 69:  members (19) 
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/sum_rename_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/sum_rename_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/root_register_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/root_register_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/base_resize_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/base_resize_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_address_resized
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_root_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_address_calculated
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_398_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	28 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/req
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(70), ack => W_fn_388_delayed_7_0_400_inst_req_0); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(28) & loadKernelChannel_CP_676_elements(72);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	76 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_update_start_
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/req
      -- 
    req_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(71), ack => W_fn_388_delayed_7_0_400_inst_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(73) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	25 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/ack
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_388_delayed_7_0_400_inst_ack_0, ack => loadKernelChannel_CP_676_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/ack
      -- 
    ack_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_388_delayed_7_0_400_inst_ack_1, ack => loadKernelChannel_CP_676_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	69 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/rr
      -- 
    rr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(74), ack => ptr_deref_406_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(73) & loadKernelChannel_CP_676_elements(69) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	21 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_update_start_
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/$entry
      -- 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(75), ack => ptr_deref_406_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(77);
      gj_loadKernelChannel_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	64 
    -- CP-element group 76: 	71 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/ra
      -- 
    ra_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	87 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	42 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/merge_ack
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/merge_req
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/$entry
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/ca
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/$exit
      -- 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	28 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/req
      -- 
    req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(78), ack => W_fn_394_delayed_13_0_408_inst_req_0); -- 
    loadKernelChannel_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(28) & loadKernelChannel_CP_676_elements(80);
      gj_loadKernelChannel_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	21 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_update_start_
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/req
      -- 
    req_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(79), ack => W_fn_394_delayed_13_0_408_inst_req_1); -- 
    loadKernelChannel_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(81);
      gj_loadKernelChannel_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	25 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/ack
      -- 
    ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_394_delayed_13_0_408_inst_ack_0, ack => loadKernelChannel_CP_676_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	87 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	42 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/ack
      -- 
    ack_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_394_delayed_13_0_408_inst_ack_1, ack => loadKernelChannel_CP_676_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	46 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/req
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/$entry
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(82), ack => W_fetch_val_396_delayed_13_0_411_inst_req_0); -- 
    loadKernelChannel_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	21 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_update_start_
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/req
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/$entry
      -- 
    req_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(83), ack => W_fetch_val_396_delayed_13_0_411_inst_req_1); -- 
    loadKernelChannel_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(85);
      gj_loadKernelChannel_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/ack
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/$exit
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_396_delayed_13_0_411_inst_ack_0, ack => loadKernelChannel_CP_676_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	42 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_update_completed_
      -- 
    ack_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_396_delayed_13_0_411_inst_ack_1, ack => loadKernelChannel_CP_676_elements(85)); -- 
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	18 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	19 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_676_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_676_elements(18), ack => loadKernelChannel_CP_676_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	21 
    -- CP-element group 87: 	77 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	62 
    -- CP-element group 87: 	81 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	15 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(62) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85);
      gj_loadKernelChannel_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	14 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/$exit
      -- CP-element group 88: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/ack
      -- 
    ack_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_350_branch_ack_0, ack => loadKernelChannel_CP_676_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	14 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/$exit
      -- CP-element group 89: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/ack
      -- 
    ack_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_350_branch_ack_1, ack => loadKernelChannel_CP_676_elements(89)); -- 
    -- CP-element group 90:  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	12 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	10 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_349/do_while_stmt_350/$exit
      -- 
    loadKernelChannel_CP_676_elements(90) <= loadKernelChannel_CP_676_elements(12);
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	10 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_Sample/ra
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_Sample/$exit
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_sample_completed_
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_0, ack => loadKernelChannel_CP_676_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	10 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_Update/$exit
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_sample_start_
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_update_completed_
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/req
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_Update/ca
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_1, ack => loadKernelChannel_CP_676_elements(92)); -- 
    req_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(92), ack => WPIPE_size_pipe_428_inst_req_0); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/ack
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_sample_completed_
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/req
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_update_start_
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/$exit
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/$entry
      -- 
    ack_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_428_inst_ack_0, ack => loadKernelChannel_CP_676_elements(93)); -- 
    req_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(93), ack => WPIPE_size_pipe_428_inst_req_1); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 assign_stmt_433/$exit
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/ack
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_update_completed_
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/$exit
      -- CP-element group 94: 	 $exit
      -- 
    ack_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_428_inst_ack_1, ack => loadKernelChannel_CP_676_elements(94)); -- 
    loadKernelChannel_do_while_stmt_350_terminator_1088: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_350_terminator_1088", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_676_elements(15),loop_continue => loadKernelChannel_CP_676_elements(89),loop_terminate => loadKernelChannel_CP_676_elements(88),loop_back => loadKernelChannel_CP_676_elements(13),loop_exit => loadKernelChannel_CP_676_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_352_phi_seq_872_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(29);
      loadKernelChannel_CP_676_elements(34)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(36);
      loadKernelChannel_CP_676_elements(35)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(37);
      loadKernelChannel_CP_676_elements(30) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(31);
      loadKernelChannel_CP_676_elements(38)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(40);
      loadKernelChannel_CP_676_elements(39)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(41);
      loadKernelChannel_CP_676_elements(32) <= phi_mux_reqs(1);
      phi_stmt_352_phi_seq_872 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_352_phi_seq_872") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(26), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(27), 
          phi_update_req => loadKernelChannel_CP_676_elements(22), 
          phi_update_ack => loadKernelChannel_CP_676_elements(28), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(33), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_356_phi_seq_926_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(47);
      loadKernelChannel_CP_676_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(54);
      loadKernelChannel_CP_676_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(55);
      loadKernelChannel_CP_676_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(49);
      loadKernelChannel_CP_676_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(58);
      loadKernelChannel_CP_676_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(59);
      loadKernelChannel_CP_676_elements(50) <= phi_mux_reqs(1);
      phi_stmt_356_phi_seq_926 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_356_phi_seq_926") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(44), 
          phi_update_req => loadKernelChannel_CP_676_elements(45), 
          phi_update_ack => loadKernelChannel_CP_676_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_814_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_676_elements(16);
        preds(1)  <= loadKernelChannel_CP_676_elements(17);
        entry_tmerge_814 : transition_merge -- 
          generic map(name => " entry_tmerge_814")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_676_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_365_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_387_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_378_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_396_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_396_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_396_wire : std_logic_vector(63 downto 0);
    signal R_sh_start_332_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_332_scaled : std_logic_vector(13 downto 0);
    signal SUB_u64_u64_366_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_424_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_431_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_425_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_333_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_root_address : std_logic_vector(13 downto 0);
    signal fetch_addr_335 : std_logic_vector(31 downto 0);
    signal fetch_addr_399 : std_logic_vector(31 downto 0);
    signal fetch_val_356 : std_logic_vector(63 downto 0);
    signal fetch_val_396_delayed_13_0_413 : std_logic_vector(63 downto 0);
    signal first_fill_344 : std_logic_vector(0 downto 0);
    signal fn_388_delayed_7_0_402 : std_logic_vector(0 downto 0);
    signal fn_390 : std_logic_vector(0 downto 0);
    signal fn_394_delayed_13_0_410 : std_logic_vector(0 downto 0);
    signal fv_407 : std_logic_vector(63 downto 0);
    signal konst_326_wire_constant : std_logic_vector(63 downto 0);
    signal konst_342_wire_constant : std_logic_vector(63 downto 0);
    signal konst_362_wire_constant : std_logic_vector(63 downto 0);
    signal konst_364_wire_constant : std_logic_vector(63 downto 0);
    signal konst_367_wire_constant : std_logic_vector(63 downto 0);
    signal konst_372_wire_constant : std_logic_vector(63 downto 0);
    signal konst_386_wire_constant : std_logic_vector(63 downto 0);
    signal konst_388_wire_constant : std_logic_vector(63 downto 0);
    signal konst_395_wire_constant : std_logic_vector(63 downto 0);
    signal konst_423_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_339 : std_logic_vector(63 downto 0);
    signal my_fetch_339_359_buffered : std_logic_vector(63 downto 0);
    signal my_num1_369 : std_logic_vector(63 downto 0);
    signal mycount_352 : std_logic_vector(63 downto 0);
    signal nfetch_val_419 : std_logic_vector(63 downto 0);
    signal nfetch_val_419_358_buffered : std_logic_vector(63 downto 0);
    signal nmycount_374 : std_logic_vector(63 downto 0);
    signal nmycount_374_354_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_338_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_338_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_338_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_338_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_338_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_406_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_406_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_406_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_406_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_406_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_start_328 : std_logic_vector(63 downto 0);
    signal start_add_355_buffered : std_logic_vector(63 downto 0);
    signal start_next_348 : std_logic_vector(0 downto 0);
    signal type_cast_432_wire : std_logic_vector(31 downto 0);
    signal var_val_380 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_333_constant_part_of_offset <= "00000000000000";
    array_obj_ref_333_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_333_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_333_resized_base_address <= "00000000000000";
    array_obj_ref_397_constant_part_of_offset <= "00000000000000";
    array_obj_ref_397_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_397_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_397_resized_base_address <= "00000000000000";
    konst_326_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_342_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_362_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_364_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_367_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_372_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_388_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_395_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_423_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_338_word_offset_0 <= "00000000000000";
    ptr_deref_406_word_offset_0 <= "00000000000000";
    phi_stmt_352: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_374_354_buffered & start_add_355_buffered;
      req <= phi_stmt_352_req_0 & phi_stmt_352_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_352",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_352_ack_0,
          idata => idata,
          odata => mycount_352,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_352
    phi_stmt_356: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_419_358_buffered & my_fetch_339_359_buffered;
      req <= phi_stmt_356_req_0 & phi_stmt_356_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_356",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_356_ack_0,
          idata => idata,
          odata => fetch_val_356,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_356
    -- flow-through select operator MUX_418_inst
    nfetch_val_419 <= fv_407 when (fn_394_delayed_13_0_410(0) /=  '0') else fetch_val_396_delayed_13_0_413;
    W_fetch_val_396_delayed_13_0_411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_396_delayed_13_0_411_inst_req_0;
      W_fetch_val_396_delayed_13_0_411_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_396_delayed_13_0_411_inst_req_1;
      W_fetch_val_396_delayed_13_0_411_inst_ack_1<= rack(0);
      W_fetch_val_396_delayed_13_0_411_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_396_delayed_13_0_411_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_396_delayed_13_0_413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_388_delayed_7_0_400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_388_delayed_7_0_400_inst_req_0;
      W_fn_388_delayed_7_0_400_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_388_delayed_7_0_400_inst_req_1;
      W_fn_388_delayed_7_0_400_inst_ack_1<= rack(0);
      W_fn_388_delayed_7_0_400_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_388_delayed_7_0_400_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_388_delayed_7_0_402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_394_delayed_13_0_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_394_delayed_13_0_408_inst_req_0;
      W_fn_394_delayed_13_0_408_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_394_delayed_13_0_408_inst_req_1;
      W_fn_394_delayed_13_0_408_inst_ack_1<= rack(0);
      W_fn_394_delayed_13_0_408_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_394_delayed_13_0_408_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_394_delayed_13_0_410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_334_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_334_final_reg_req_0;
      addr_of_334_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_334_final_reg_req_1;
      addr_of_334_final_reg_ack_1<= rack(0);
      addr_of_334_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_334_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_333_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_335,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_398_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_398_final_reg_req_0;
      addr_of_398_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_398_final_reg_req_1;
      addr_of_398_final_reg_ack_1<= rack(0);
      addr_of_398_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_398_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_397_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_339_359_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_339_359_buf_req_0;
      my_fetch_339_359_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_339_359_buf_req_1;
      my_fetch_339_359_buf_ack_1<= rack(0);
      my_fetch_339_359_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_339_359_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_339_359_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_419_358_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_419_358_buf_req_0;
      nfetch_val_419_358_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_419_358_buf_req_1;
      nfetch_val_419_358_buf_ack_1<= rack(0);
      nfetch_val_419_358_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_419_358_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_419_358_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_374_354_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_374_354_buf_req_0;
      nmycount_374_354_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_374_354_buf_req_1;
      nmycount_374_354_buf_ack_1<= rack(0);
      nmycount_374_354_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_374_354_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_374_354_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_355_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_355_buf_req_0;
      start_add_355_buf_ack_0<= wack(0);
      rreq(0) <= start_add_355_buf_req_1;
      start_add_355_buf_ack_1<= rack(0);
      start_add_355_buf : InterlockBuffer generic map ( -- 
        name => "start_add_355_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_355_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_379_inst
    process(LSHR_u64_u64_378_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_378_wire(15 downto 0);
      var_val_380 <= tmp_var; -- 
    end process;
    type_cast_432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_432_inst_req_0;
      type_cast_432_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_432_inst_req_1;
      type_cast_432_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  first_fill_344(0);
      type_cast_432_inst_gI: SplitGuardInterface generic map(name => "type_cast_432_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SUB_u64_u64_431_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_432_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_333_index_1_rename
    process(R_sh_start_332_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_332_resized;
      ov(13 downto 0) := iv;
      R_sh_start_332_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_333_index_1_resize
    process(sh_start_328) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_328;
      ov := iv(13 downto 0);
      R_sh_start_332_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_333_root_address_inst
    process(array_obj_ref_333_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_333_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_333_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_index_1_rename
    process(LSHR_u64_u64_396_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_396_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_396_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_index_1_resize
    process(LSHR_u64_u64_396_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_396_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_396_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_root_address_inst
    process(array_obj_ref_397_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_397_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_397_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_addr_0
    process(ptr_deref_338_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_338_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_base_resize
    process(fetch_addr_335) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_335;
      ov := iv(13 downto 0);
      ptr_deref_338_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_gather_scatter
    process(ptr_deref_338_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_data_0;
      ov(63 downto 0) := iv;
      my_fetch_339 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_root_address_inst
    process(ptr_deref_338_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_338_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_addr_0
    process(ptr_deref_406_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_406_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_base_resize
    process(fetch_addr_399) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_399;
      ov := iv(13 downto 0);
      ptr_deref_406_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_gather_scatter
    process(ptr_deref_406_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_data_0;
      ov(63 downto 0) := iv;
      fv_407 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_root_address_inst
    process(ptr_deref_406_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_406_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_350_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_425_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_350_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_350_branch_req_0,
          ack0 => do_while_stmt_350_branch_ack_0,
          ack1 => do_while_stmt_350_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_373_inst
    process(mycount_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_352, konst_372_wire_constant, tmp_var);
      nmycount_374 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_365_inst
    process(mycount_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_352, konst_364_wire_constant, tmp_var);
      AND_u64_u64_365_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_387_inst
    process(nmycount_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_374, konst_386_wire_constant, tmp_var);
      AND_u64_u64_387_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_343_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_342_wire_constant, tmp_var);
      first_fill_344 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_389_inst
    process(AND_u64_u64_387_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_387_wire, konst_388_wire_constant, tmp_var);
      fn_390 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_327_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_326_wire_constant, tmp_var);
      sh_start_328 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_378_inst
    process(fetch_val_356, my_num1_369) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_356, my_num1_369, tmp_var);
      LSHR_u64_u64_378_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_396_inst
    process(nmycount_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_374, konst_395_wire_constant, tmp_var);
      LSHR_u64_u64_396_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_368_inst
    process(SUB_u64_u64_366_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_366_wire, konst_367_wire_constant, tmp_var);
      my_num1_369 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_366_inst
    process(konst_362_wire_constant, AND_u64_u64_365_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_362_wire_constant, AND_u64_u64_365_wire, tmp_var);
      SUB_u64_u64_366_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_424_inst
    process(end_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, konst_423_wire_constant, tmp_var);
      SUB_u64_u64_424_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_431_inst
    process(end_add_buffer, start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, start_add_buffer, tmp_var);
      SUB_u64_u64_431_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_425_inst
    process(mycount_352, SUB_u64_u64_424_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_352, SUB_u64_u64_424_wire, tmp_var);
      ULT_u64_u1_425_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : array_obj_ref_333_index_offset 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_332_scaled;
      array_obj_ref_333_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_333_index_offset_req_0;
      array_obj_ref_333_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_333_index_offset_req_1;
      array_obj_ref_333_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_397_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_396_scaled;
      array_obj_ref_397_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_397_index_offset_req_0;
      array_obj_ref_397_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_397_index_offset_req_1;
      array_obj_ref_397_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_338_load_0 ptr_deref_406_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_338_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_406_load_0_req_0;
      ptr_deref_338_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_406_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_338_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_406_load_0_req_1;
      ptr_deref_338_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_406_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_388_delayed_7_0_402(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_338_word_address_0 & ptr_deref_406_word_address_0;
      ptr_deref_338_data_0 <= data_out(127 downto 64);
      ptr_deref_406_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_347_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_347_inst_req_0;
      RPIPE_input_done_pipe_347_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_347_inst_req_1;
      RPIPE_input_done_pipe_347_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_344(0);
      start_next_348 <= data_out(0 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_381_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_381_inst_req_0;
      WPIPE_kernel_pipe1_381_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_381_inst_req_1;
      WPIPE_kernel_pipe1_381_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val_380;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_size_pipe_428_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_428_inst_req_0;
      WPIPE_size_pipe_428_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_428_inst_req_1;
      WPIPE_size_pipe_428_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= first_fill_344(0);
      data_in <= type_cast_432_wire;
      size_pipe_write_1_gI: SplitGuardInterface generic map(name => "size_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_637_start: Boolean;
  signal timer_CP_637_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_318_load_0_req_0 : boolean;
  signal LOAD_count_318_load_0_ack_0 : boolean;
  signal LOAD_count_318_load_0_req_1 : boolean;
  signal LOAD_count_318_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_637_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_637: Block -- control-path 
    signal timer_CP_637_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_637_elements(0) <= timer_CP_637_start;
    timer_CP_637_symbol <= timer_CP_637_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_319/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_sample_start_
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_update_start_
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/cr
      -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_318_load_0_req_1); -- 
    rr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_318_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_sample_completed_
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/ra
      -- 
    ra_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_318_load_0_ack_0, ack => timer_CP_637_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_319/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_update_completed_
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/merge_ack
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_318_load_0_ack_1, ack => timer_CP_637_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_318_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_318_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_318_word_address_0 <= "0";
    -- equivalence LOAD_count_318_gather_scatter
    process(LOAD_count_318_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_318_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_318_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_318_load_0_req_0;
      LOAD_count_318_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_318_load_0_req_1;
      LOAD_count_318_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_318_word_address_0;
      LOAD_count_318_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_5094_start: Boolean;
  signal timerDaemon_CP_5094_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_2114_branch_req_0 : boolean;
  signal phi_stmt_2116_req_1 : boolean;
  signal phi_stmt_2116_req_0 : boolean;
  signal phi_stmt_2116_ack_0 : boolean;
  signal ADD_u64_u64_2122_inst_req_0 : boolean;
  signal ADD_u64_u64_2122_inst_ack_0 : boolean;
  signal ADD_u64_u64_2122_inst_req_1 : boolean;
  signal ADD_u64_u64_2122_inst_ack_1 : boolean;
  signal STORE_count_2124_store_0_req_0 : boolean;
  signal STORE_count_2124_store_0_ack_0 : boolean;
  signal STORE_count_2124_store_0_req_1 : boolean;
  signal STORE_count_2124_store_0_ack_1 : boolean;
  signal do_while_stmt_2114_branch_ack_0 : boolean;
  signal do_while_stmt_2114_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_5094_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_5094_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_5094_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_5094_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_5094: Block -- control-path 
    signal timerDaemon_CP_5094_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_5094_elements(0) <= timerDaemon_CP_5094_start;
    timerDaemon_CP_5094_symbol <= timerDaemon_CP_5094_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2113/$entry
      -- CP-element group 0: 	 branch_block_stmt_2113/branch_block_stmt_2113__entry__
      -- CP-element group 0: 	 branch_block_stmt_2113/do_while_stmt_2114__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2113/$exit
      -- CP-element group 1: 	 branch_block_stmt_2113/branch_block_stmt_2113__exit__
      -- CP-element group 1: 	 branch_block_stmt_2113/do_while_stmt_2114__exit__
      -- 
    timerDaemon_CP_5094_elements(1) <= timerDaemon_CP_5094_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2113/do_while_stmt_2114/$entry
      -- CP-element group 2: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114__entry__
      -- 
    timerDaemon_CP_5094_elements(2) <= timerDaemon_CP_5094_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114__exit__
      -- 
    -- Element group timerDaemon_CP_5094_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2113/do_while_stmt_2114/loop_back
      -- 
    -- Element group timerDaemon_CP_5094_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2113/do_while_stmt_2114/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2113/do_while_stmt_2114/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2113/do_while_stmt_2114/loop_taken/$entry
      -- 
    timerDaemon_CP_5094_elements(5) <= timerDaemon_CP_5094_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2113/do_while_stmt_2114/loop_body_done
      -- 
    timerDaemon_CP_5094_elements(6) <= timerDaemon_CP_5094_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_5094_elements(7) <= timerDaemon_CP_5094_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_5094_elements(8) <= timerDaemon_CP_5094_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	31 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_5094_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	35 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/condition_evaluated
      -- 
    condition_evaluated_5118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_5118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5094_elements(10), ack => do_while_stmt_2114_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5094_elements(15) & timerDaemon_CP_5094_elements(35);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5094_elements(12) & timerDaemon_CP_5094_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5094_elements(9) & timerDaemon_CP_5094_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_update_start_
      -- CP-element group 13: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5094_elements(9) & timerDaemon_CP_5094_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_5094_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_5094_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_loopback_trigger
      -- 
    timerDaemon_CP_5094_elements(16) <= timerDaemon_CP_5094_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_loopback_sample_req_ps
      -- 
    phi_stmt_2116_loopback_sample_req_5133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2116_loopback_sample_req_5133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5094_elements(17), ack => phi_stmt_2116_req_1); -- 
    -- Element group timerDaemon_CP_5094_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_entry_trigger
      -- 
    timerDaemon_CP_5094_elements(18) <= timerDaemon_CP_5094_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_entry_sample_req_ps
      -- 
    phi_stmt_2116_entry_sample_req_5136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2116_entry_sample_req_5136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5094_elements(19), ack => phi_stmt_2116_req_0); -- 
    -- Element group timerDaemon_CP_5094_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/phi_stmt_2116_phi_mux_ack_ps
      -- 
    phi_stmt_2116_phi_mux_ack_5139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2116_ack_0, ack => timerDaemon_CP_5094_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/type_cast_2119_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/type_cast_2119_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/type_cast_2119_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/type_cast_2119_sample_completed_
      -- 
    -- Element group timerDaemon_CP_5094_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/type_cast_2119_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/type_cast_2119_update_start_
      -- 
    -- Element group timerDaemon_CP_5094_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/type_cast_2119_update_completed__ps
      -- 
    timerDaemon_CP_5094_elements(23) <= timerDaemon_CP_5094_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/type_cast_2119_update_completed_
      -- 
    -- Element group timerDaemon_CP_5094_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_5094_elements(22), ack => timerDaemon_CP_5094_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_5094_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_update_start__ps
      -- 
    -- Element group timerDaemon_CP_5094_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_Sample/rr
      -- 
    rr_5160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5094_elements(27), ack => ADD_u64_u64_2122_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5094_elements(25) & timerDaemon_CP_5094_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_Update/cr
      -- 
    cr_5165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5094_elements(28), ack => ADD_u64_u64_2122_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5094_elements(26) & timerDaemon_CP_5094_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_Sample/ra
      -- 
    ra_5161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2122_inst_ack_0, ack => timerDaemon_CP_5094_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/ADD_u64_u64_2122_Update/ca
      -- 
    ca_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2122_inst_ack_1, ack => timerDaemon_CP_5094_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/STORE_count_2124_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/STORE_count_2124_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/STORE_count_2124_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/STORE_count_2124_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/word_access_start/word_0/rr
      -- 
    rr_5188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5094_elements(31), ack => STORE_count_2124_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_5094_elements(9) & timerDaemon_CP_5094_elements(15) & timerDaemon_CP_5094_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Update/word_access_complete/word_0/cr
      -- 
    cr_5199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5094_elements(32), ack => STORE_count_2124_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_5094_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Sample/word_access_start/word_0/ra
      -- 
    ra_5189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2124_store_0_ack_0, ack => timerDaemon_CP_5094_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/STORE_count_2124_Update/word_access_complete/word_0/ca
      -- 
    ca_5200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2124_store_0_ack_1, ack => timerDaemon_CP_5094_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_5094_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_5094_elements(9), ack => timerDaemon_CP_5094_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_2113/do_while_stmt_2114/do_while_stmt_2114_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5094_elements(14) & timerDaemon_CP_5094_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5094_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_2113/do_while_stmt_2114/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_2113/do_while_stmt_2114/loop_exit/ack
      -- 
    ack_5205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2114_branch_ack_0, ack => timerDaemon_CP_5094_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_2113/do_while_stmt_2114/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_2113/do_while_stmt_2114/loop_taken/ack
      -- 
    ack_5209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2114_branch_ack_1, ack => timerDaemon_CP_5094_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2113/do_while_stmt_2114/$exit
      -- 
    timerDaemon_CP_5094_elements(39) <= timerDaemon_CP_5094_elements(3);
    timerDaemon_do_while_stmt_2114_terminator_5210: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2114_terminator_5210", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_5094_elements(6),loop_continue => timerDaemon_CP_5094_elements(38),loop_terminate => timerDaemon_CP_5094_elements(37),loop_back => timerDaemon_CP_5094_elements(4),loop_exit => timerDaemon_CP_5094_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2116_phi_seq_5167_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_5094_elements(18);
      timerDaemon_CP_5094_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_5094_elements(21);
      timerDaemon_CP_5094_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_5094_elements(23);
      timerDaemon_CP_5094_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_5094_elements(16);
      timerDaemon_CP_5094_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_5094_elements(29);
      timerDaemon_CP_5094_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_5094_elements(30);
      timerDaemon_CP_5094_elements(17) <= phi_mux_reqs(1);
      phi_stmt_2116_phi_seq_5167 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_2116_phi_seq_5167") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_5094_elements(11), 
          phi_sample_ack => timerDaemon_CP_5094_elements(14), 
          phi_update_req => timerDaemon_CP_5094_elements(13), 
          phi_update_ack => timerDaemon_CP_5094_elements(15), 
          phi_mux_ack => timerDaemon_CP_5094_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_5119_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_5094_elements(7);
        preds(1)  <= timerDaemon_CP_5094_elements(8);
        entry_tmerge_5119 : transition_merge -- 
          generic map(name => " entry_tmerge_5119")
          port map (preds => preds, symbol_out => timerDaemon_CP_5094_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_2122_wire : std_logic_vector(63 downto 0);
    signal STORE_count_2124_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_2124_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_2121_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2128_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_2116 : std_logic_vector(63 downto 0);
    signal type_cast_2119_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_2124_word_address_0 <= "0";
    konst_2121_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2128_wire_constant <= "1";
    type_cast_2119_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2116: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2119_wire_constant & ADD_u64_u64_2122_wire;
      req <= phi_stmt_2116_req_0 & phi_stmt_2116_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2116",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2116_ack_0,
          idata => idata,
          odata => ncount_2116,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2116
    -- equivalence STORE_count_2124_gather_scatter
    process(ncount_2116) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_2116;
      ov(63 downto 0) := iv;
      STORE_count_2124_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_2114_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2128_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2114_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2114_branch_req_0,
          ack0 => do_while_stmt_2114_branch_ack_0,
          ack1 => do_while_stmt_2114_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_2122_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_2116;
      ADD_u64_u64_2122_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2122_inst_req_0;
      ADD_u64_u64_2122_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2122_inst_req_1;
      ADD_u64_u64_2122_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_2124_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_2124_store_0_req_0;
      STORE_count_2124_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_2124_store_0_req_1;
      STORE_count_2124_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_2124_word_address_0;
      data_in <= STORE_count_2124_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_num_cont :  std_logic_vector(15 downto 0);
  signal access_T_row1 :  std_logic_vector(15 downto 0);
  signal access_T_col1 :  std_logic_vector(15 downto 0);
  signal access_T_rk1 :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(95 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(95 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(95 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_end_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(127 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(127 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_num_cont <= access_T_in_args(95 downto 80);
  access_T_row1 <= access_T_in_args(79 downto 64);
  access_T_col1 <= access_T_in_args(63 downto 48);
  access_T_rk1 <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      num_cont => access_T_num_cont,
      row1 => access_T_row1,
      col1 => access_T_col1,
      rk1 => access_T_rk1,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(95 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(127 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(31 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(0 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(127 downto 64);
  loadKernelChannel_end_add <= loadKernelChannel_in_args(63 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 128,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      end_add => loadKernelChannel_end_add,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(0 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(31 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(1 downto 1),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(1 downto 1),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(31 downto 16),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
